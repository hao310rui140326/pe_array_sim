// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Internal Build 259 12/02/2018 SJ Pro Edition"

// DATE "12/08/2018 22:19:14"

// 
// Device: Altera 10AX115S2F45I1SG Package FBGA1932
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module pe_dot_alm_a10_12x12x16 (
	dout,
	clk,
	din_a,
	din_b);
output 	[26:0] dout;
input 	clk;
input 	[191:0] din_a;
input 	[191:0] din_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire Xd_0__inst_inst_inst_rtl_1_sumout ;
wire Xd_0__inst_inst_inst_rtl_2 ;
wire Xd_0__inst_inst_inst_rtl_3 ;
wire Xd_0__inst_inst_inst_rtl_5_sumout ;
wire Xd_0__inst_inst_inst_rtl_6 ;
wire Xd_0__inst_inst_inst_rtl_7 ;
wire Xd_0__inst_inst_inst_rtl_9_sumout ;
wire Xd_0__inst_inst_inst_rtl_10 ;
wire Xd_0__inst_inst_inst_rtl_11 ;
wire Xd_0__inst_inst_inst_rtl_13_sumout ;
wire Xd_0__inst_inst_inst_rtl_14 ;
wire Xd_0__inst_inst_inst_rtl_15 ;
wire Xd_0__inst_inst_inst_rtl_17_sumout ;
wire Xd_0__inst_inst_inst_rtl_18 ;
wire Xd_0__inst_inst_inst_rtl_19 ;
wire Xd_0__inst_inst_inst_rtl_21_sumout ;
wire Xd_0__inst_inst_inst_rtl_22 ;
wire Xd_0__inst_inst_inst_rtl_23 ;
wire Xd_0__inst_inst_inst_rtl_25_sumout ;
wire Xd_0__inst_inst_inst_rtl_26 ;
wire Xd_0__inst_inst_inst_rtl_27 ;
wire Xd_0__inst_inst_inst_rtl_29_sumout ;
wire Xd_0__inst_inst_inst_rtl_30 ;
wire Xd_0__inst_inst_inst_rtl_31 ;
wire Xd_0__inst_inst_inst_rtl_33_sumout ;
wire Xd_0__inst_inst_inst_rtl_34 ;
wire Xd_0__inst_inst_inst_rtl_35 ;
wire Xd_0__inst_inst_inst_rtl_37_sumout ;
wire Xd_0__inst_inst_inst_rtl_38 ;
wire Xd_0__inst_inst_inst_rtl_39 ;
wire Xd_0__inst_inst_inst_rtl_41_sumout ;
wire Xd_0__inst_inst_inst_rtl_42 ;
wire Xd_0__inst_inst_inst_rtl_43 ;
wire Xd_0__inst_inst_inst_rtl_45_sumout ;
wire Xd_0__inst_inst_inst_rtl_46 ;
wire Xd_0__inst_inst_inst_rtl_47 ;
wire Xd_0__inst_inst_inst_rtl_49_sumout ;
wire Xd_0__inst_inst_inst_rtl_50 ;
wire Xd_0__inst_inst_inst_rtl_51 ;
wire Xd_0__inst_inst_inst_rtl_53_sumout ;
wire Xd_0__inst_inst_inst_rtl_54 ;
wire Xd_0__inst_inst_inst_rtl_55 ;
wire Xd_0__inst_inst_inst_rtl_57_sumout ;
wire Xd_0__inst_inst_inst_rtl_58 ;
wire Xd_0__inst_inst_inst_rtl_59 ;
wire Xd_0__inst_inst_inst_rtl_61_sumout ;
wire Xd_0__inst_inst_inst_rtl_62 ;
wire Xd_0__inst_inst_inst_rtl_63 ;
wire Xd_0__inst_inst_inst_rtl_65_sumout ;
wire Xd_0__inst_inst_inst_rtl_66 ;
wire Xd_0__inst_inst_inst_rtl_67 ;
wire Xd_0__inst_inst_inst_rtl_69_sumout ;
wire Xd_0__inst_inst_inst_rtl_70 ;
wire Xd_0__inst_inst_inst_rtl_71 ;
wire Xd_0__inst_inst_inst_rtl_73_sumout ;
wire Xd_0__inst_inst_inst_rtl_74 ;
wire Xd_0__inst_inst_inst_rtl_75 ;
wire Xd_0__inst_inst_inst_rtl_77_sumout ;
wire Xd_0__inst_inst_inst_rtl_78 ;
wire Xd_0__inst_inst_inst_rtl_79 ;
wire Xd_0__inst_inst_inst_rtl_81_sumout ;
wire Xd_0__inst_inst_inst_rtl_82 ;
wire Xd_0__inst_inst_inst_rtl_83 ;
wire Xd_0__inst_inst_inst_rtl_85_sumout ;
wire Xd_0__inst_inst_inst_rtl_86 ;
wire Xd_0__inst_inst_inst_rtl_87 ;
wire Xd_0__inst_inst_inst_rtl_89_sumout ;
wire Xd_0__inst_inst_inst_rtl_90 ;
wire Xd_0__inst_inst_inst_rtl_91 ;
wire Xd_0__inst_inst_inst_rtl_93_sumout ;
wire Xd_0__inst_inst_inst_rtl_94 ;
wire Xd_0__inst_inst_inst_rtl_95 ;
wire Xd_0__inst_inst_inst_rtl_97_sumout ;
wire Xd_0__inst_inst_inst_rtl_98 ;
wire Xd_0__inst_inst_inst_rtl_99 ;
wire Xd_0__inst_inst_inst_rtl_101_sumout ;
wire Xd_0__inst_inst_inst_rtl_102 ;
wire Xd_0__inst_inst_inst_rtl_103 ;
wire Xd_0__inst_inst_inst_rtl_105_sumout ;
wire Xd_0__inst_mult_4_173 ;
wire Xd_0__inst_mult_4_174 ;
wire Xd_0__inst_mult_4_175 ;
wire Xd_0__inst_inst_add_4_1_sumout ;
wire Xd_0__inst_inst_add_4_2 ;
wire Xd_0__inst_inst_add_4_3 ;
wire Xd_0__inst_inst_add_2_1_sumout ;
wire Xd_0__inst_inst_add_2_2 ;
wire Xd_0__inst_inst_add_2_3 ;
wire Xd_0__inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_add_0_2 ;
wire Xd_0__inst_inst_add_0_3 ;
wire Xd_0__inst_mult_4_177 ;
wire Xd_0__inst_mult_4_178 ;
wire Xd_0__inst_mult_4_179 ;
wire Xd_0__inst_inst_add_4_5_sumout ;
wire Xd_0__inst_inst_add_4_6 ;
wire Xd_0__inst_inst_add_4_7 ;
wire Xd_0__inst_inst_add_2_5_sumout ;
wire Xd_0__inst_inst_add_2_6 ;
wire Xd_0__inst_inst_add_2_7 ;
wire Xd_0__inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_add_0_6 ;
wire Xd_0__inst_inst_add_0_7 ;
wire Xd_0__inst_inst_add_4_9_sumout ;
wire Xd_0__inst_inst_add_4_10 ;
wire Xd_0__inst_inst_add_4_11 ;
wire Xd_0__inst_inst_add_2_9_sumout ;
wire Xd_0__inst_inst_add_2_10 ;
wire Xd_0__inst_inst_add_2_11 ;
wire Xd_0__inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_add_0_10 ;
wire Xd_0__inst_inst_add_0_11 ;
wire Xd_0__inst_inst_add_4_13_sumout ;
wire Xd_0__inst_inst_add_4_14 ;
wire Xd_0__inst_inst_add_4_15 ;
wire Xd_0__inst_inst_add_2_13_sumout ;
wire Xd_0__inst_inst_add_2_14 ;
wire Xd_0__inst_inst_add_2_15 ;
wire Xd_0__inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_add_0_14 ;
wire Xd_0__inst_inst_add_0_15 ;
wire Xd_0__inst_inst_add_4_17_sumout ;
wire Xd_0__inst_inst_add_4_18 ;
wire Xd_0__inst_inst_add_4_19 ;
wire Xd_0__inst_inst_add_2_17_sumout ;
wire Xd_0__inst_inst_add_2_18 ;
wire Xd_0__inst_inst_add_2_19 ;
wire Xd_0__inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_add_0_18 ;
wire Xd_0__inst_inst_add_0_19 ;
wire Xd_0__inst_inst_add_4_21_sumout ;
wire Xd_0__inst_inst_add_4_22 ;
wire Xd_0__inst_inst_add_4_23 ;
wire Xd_0__inst_inst_add_2_21_sumout ;
wire Xd_0__inst_inst_add_2_22 ;
wire Xd_0__inst_inst_add_2_23 ;
wire Xd_0__inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_add_0_22 ;
wire Xd_0__inst_inst_add_0_23 ;
wire Xd_0__inst_inst_add_4_25_sumout ;
wire Xd_0__inst_inst_add_4_26 ;
wire Xd_0__inst_inst_add_4_27 ;
wire Xd_0__inst_inst_add_2_25_sumout ;
wire Xd_0__inst_inst_add_2_26 ;
wire Xd_0__inst_inst_add_2_27 ;
wire Xd_0__inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_add_0_26 ;
wire Xd_0__inst_inst_add_0_27 ;
wire Xd_0__inst_inst_add_4_29_sumout ;
wire Xd_0__inst_inst_add_4_30 ;
wire Xd_0__inst_inst_add_4_31 ;
wire Xd_0__inst_inst_add_2_29_sumout ;
wire Xd_0__inst_inst_add_2_30 ;
wire Xd_0__inst_inst_add_2_31 ;
wire Xd_0__inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_add_0_30 ;
wire Xd_0__inst_inst_add_0_31 ;
wire Xd_0__inst_inst_add_4_33_sumout ;
wire Xd_0__inst_inst_add_4_34 ;
wire Xd_0__inst_inst_add_4_35 ;
wire Xd_0__inst_inst_add_2_33_sumout ;
wire Xd_0__inst_inst_add_2_34 ;
wire Xd_0__inst_inst_add_2_35 ;
wire Xd_0__inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_add_0_34 ;
wire Xd_0__inst_inst_add_0_35 ;
wire Xd_0__inst_inst_add_4_37_sumout ;
wire Xd_0__inst_inst_add_4_38 ;
wire Xd_0__inst_inst_add_4_39 ;
wire Xd_0__inst_inst_add_2_37_sumout ;
wire Xd_0__inst_inst_add_2_38 ;
wire Xd_0__inst_inst_add_2_39 ;
wire Xd_0__inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_add_0_38 ;
wire Xd_0__inst_inst_add_0_39 ;
wire Xd_0__inst_inst_add_4_41_sumout ;
wire Xd_0__inst_inst_add_4_42 ;
wire Xd_0__inst_inst_add_4_43 ;
wire Xd_0__inst_inst_add_2_41_sumout ;
wire Xd_0__inst_inst_add_2_42 ;
wire Xd_0__inst_inst_add_2_43 ;
wire Xd_0__inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_add_0_42 ;
wire Xd_0__inst_inst_add_0_43 ;
wire Xd_0__inst_inst_add_4_45_sumout ;
wire Xd_0__inst_inst_add_4_46 ;
wire Xd_0__inst_inst_add_4_47 ;
wire Xd_0__inst_inst_add_2_45_sumout ;
wire Xd_0__inst_inst_add_2_46 ;
wire Xd_0__inst_inst_add_2_47 ;
wire Xd_0__inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_add_0_46 ;
wire Xd_0__inst_inst_add_0_47 ;
wire Xd_0__inst_inst_add_4_49_sumout ;
wire Xd_0__inst_inst_add_4_50 ;
wire Xd_0__inst_inst_add_4_51 ;
wire Xd_0__inst_inst_add_2_49_sumout ;
wire Xd_0__inst_inst_add_2_50 ;
wire Xd_0__inst_inst_add_2_51 ;
wire Xd_0__inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_add_0_50 ;
wire Xd_0__inst_inst_add_0_51 ;
wire Xd_0__inst_inst_add_4_53_sumout ;
wire Xd_0__inst_inst_add_4_54 ;
wire Xd_0__inst_inst_add_4_55 ;
wire Xd_0__inst_inst_add_2_53_sumout ;
wire Xd_0__inst_inst_add_2_54 ;
wire Xd_0__inst_inst_add_2_55 ;
wire Xd_0__inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_add_0_54 ;
wire Xd_0__inst_inst_add_0_55 ;
wire Xd_0__inst_inst_add_4_57_sumout ;
wire Xd_0__inst_inst_add_4_58 ;
wire Xd_0__inst_inst_add_4_59 ;
wire Xd_0__inst_inst_add_2_57_sumout ;
wire Xd_0__inst_inst_add_2_58 ;
wire Xd_0__inst_inst_add_2_59 ;
wire Xd_0__inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_add_0_58 ;
wire Xd_0__inst_inst_add_0_59 ;
wire Xd_0__inst_inst_add_4_61_sumout ;
wire Xd_0__inst_inst_add_4_62 ;
wire Xd_0__inst_inst_add_4_63 ;
wire Xd_0__inst_inst_add_2_61_sumout ;
wire Xd_0__inst_inst_add_2_62 ;
wire Xd_0__inst_inst_add_2_63 ;
wire Xd_0__inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_add_0_62 ;
wire Xd_0__inst_inst_add_0_63 ;
wire Xd_0__inst_inst_add_4_65_sumout ;
wire Xd_0__inst_inst_add_4_66 ;
wire Xd_0__inst_inst_add_4_67 ;
wire Xd_0__inst_inst_add_2_65_sumout ;
wire Xd_0__inst_inst_add_2_66 ;
wire Xd_0__inst_inst_add_2_67 ;
wire Xd_0__inst_inst_add_0_65_sumout ;
wire Xd_0__inst_inst_add_0_66 ;
wire Xd_0__inst_inst_add_0_67 ;
wire Xd_0__inst_inst_add_4_69_sumout ;
wire Xd_0__inst_inst_add_4_70 ;
wire Xd_0__inst_inst_add_4_71 ;
wire Xd_0__inst_inst_add_2_69_sumout ;
wire Xd_0__inst_inst_add_2_70 ;
wire Xd_0__inst_inst_add_2_71 ;
wire Xd_0__inst_inst_add_0_69_sumout ;
wire Xd_0__inst_inst_add_0_70 ;
wire Xd_0__inst_inst_add_0_71 ;
wire Xd_0__inst_inst_add_4_73_sumout ;
wire Xd_0__inst_inst_add_4_74 ;
wire Xd_0__inst_inst_add_4_75 ;
wire Xd_0__inst_inst_add_2_73_sumout ;
wire Xd_0__inst_inst_add_2_74 ;
wire Xd_0__inst_inst_add_2_75 ;
wire Xd_0__inst_inst_add_0_73_sumout ;
wire Xd_0__inst_inst_add_0_74 ;
wire Xd_0__inst_inst_add_0_75 ;
wire Xd_0__inst_inst_add_4_77_sumout ;
wire Xd_0__inst_inst_add_4_78 ;
wire Xd_0__inst_inst_add_4_79 ;
wire Xd_0__inst_inst_add_2_77_sumout ;
wire Xd_0__inst_inst_add_2_78 ;
wire Xd_0__inst_inst_add_2_79 ;
wire Xd_0__inst_inst_add_0_77_sumout ;
wire Xd_0__inst_inst_add_0_78 ;
wire Xd_0__inst_inst_add_0_79 ;
wire Xd_0__inst_inst_add_4_81_sumout ;
wire Xd_0__inst_inst_add_4_82 ;
wire Xd_0__inst_inst_add_4_83 ;
wire Xd_0__inst_inst_add_2_81_sumout ;
wire Xd_0__inst_inst_add_2_82 ;
wire Xd_0__inst_inst_add_2_83 ;
wire Xd_0__inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_add_0_82 ;
wire Xd_0__inst_inst_add_0_83 ;
wire Xd_0__inst_inst_add_4_85_sumout ;
wire Xd_0__inst_inst_add_4_86 ;
wire Xd_0__inst_inst_add_4_87 ;
wire Xd_0__inst_inst_add_2_85_sumout ;
wire Xd_0__inst_inst_add_2_86 ;
wire Xd_0__inst_inst_add_2_87 ;
wire Xd_0__inst_inst_add_0_85_sumout ;
wire Xd_0__inst_inst_add_0_86 ;
wire Xd_0__inst_inst_add_0_87 ;
wire Xd_0__inst_inst_add_4_89_sumout ;
wire Xd_0__inst_inst_add_4_90 ;
wire Xd_0__inst_inst_add_4_91 ;
wire Xd_0__inst_inst_add_2_89_sumout ;
wire Xd_0__inst_inst_add_2_90 ;
wire Xd_0__inst_inst_add_2_91 ;
wire Xd_0__inst_inst_add_0_89_sumout ;
wire Xd_0__inst_inst_add_0_90 ;
wire Xd_0__inst_inst_add_0_91 ;
wire Xd_0__inst_inst_add_4_93_sumout ;
wire Xd_0__inst_inst_add_4_94 ;
wire Xd_0__inst_inst_add_4_95 ;
wire Xd_0__inst_inst_add_2_93_sumout ;
wire Xd_0__inst_inst_add_2_94 ;
wire Xd_0__inst_inst_add_2_95 ;
wire Xd_0__inst_inst_add_0_93_sumout ;
wire Xd_0__inst_inst_add_0_94 ;
wire Xd_0__inst_inst_add_0_95 ;
wire Xd_0__inst_inst_add_4_97_sumout ;
wire Xd_0__inst_inst_add_2_97_sumout ;
wire Xd_0__inst_inst_add_2_98 ;
wire Xd_0__inst_inst_add_2_99 ;
wire Xd_0__inst_inst_add_0_97_sumout ;
wire Xd_0__inst_inst_add_0_98 ;
wire Xd_0__inst_inst_add_0_99 ;
wire Xd_0__inst_inst_add_2_101_sumout ;
wire Xd_0__inst_inst_add_0_101_sumout ;
wire Xd_0__inst_mult_14_173 ;
wire Xd_0__inst_mult_14_174 ;
wire Xd_0__inst_mult_14_175 ;
wire Xd_0__inst_mult_15_173 ;
wire Xd_0__inst_mult_15_174 ;
wire Xd_0__inst_mult_15_175 ;
wire Xd_0__inst_mult_12_169 ;
wire Xd_0__inst_mult_12_170 ;
wire Xd_0__inst_mult_12_171 ;
wire Xd_0__inst_mult_4_180 ;
wire Xd_0__inst_mult_4_181 ;
wire Xd_0__inst_mult_4_182 ;
wire Xd_0__inst_a1_6__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_14_177 ;
wire Xd_0__inst_mult_14_178 ;
wire Xd_0__inst_mult_14_179 ;
wire Xd_0__inst_a1_5__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_15_177 ;
wire Xd_0__inst_mult_15_178 ;
wire Xd_0__inst_mult_15_179 ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_12_173 ;
wire Xd_0__inst_mult_12_174 ;
wire Xd_0__inst_mult_12_175 ;
wire Xd_0__inst_mult_4_184 ;
wire Xd_0__inst_mult_4_185 ;
wire Xd_0__inst_mult_4_186 ;
wire Xd_0__inst_a1_6__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_mult_9_169 ;
wire Xd_0__inst_mult_9_170 ;
wire Xd_0__inst_mult_9_171 ;
wire Xd_0__inst_mult_6_169 ;
wire Xd_0__inst_mult_6_170 ;
wire Xd_0__inst_mult_6_171 ;
wire Xd_0__inst_mult_14_180 ;
wire Xd_0__inst_mult_14_184 ;
wire Xd_0__inst_mult_14_185 ;
wire Xd_0__inst_mult_14_186 ;
wire Xd_0__inst_mult_8_173 ;
wire Xd_0__inst_mult_8_174 ;
wire Xd_0__inst_mult_8_175 ;
wire Xd_0__inst_mult_11_173 ;
wire Xd_0__inst_mult_11_174 ;
wire Xd_0__inst_mult_11_175 ;
wire Xd_0__inst_mult_10_169 ;
wire Xd_0__inst_mult_10_170 ;
wire Xd_0__inst_mult_10_171 ;
wire Xd_0__inst_mult_15_180 ;
wire Xd_0__inst_mult_15_181 ;
wire Xd_0__inst_mult_15_182 ;
wire Xd_0__inst_mult_13_173 ;
wire Xd_0__inst_mult_13_174 ;
wire Xd_0__inst_mult_13_175 ;
wire Xd_0__inst_mult_15_184 ;
wire Xd_0__inst_mult_15_185 ;
wire Xd_0__inst_mult_15_186 ;
wire Xd_0__inst_mult_12_176 ;
wire Xd_0__inst_mult_12_177 ;
wire Xd_0__inst_mult_12_178 ;
wire Xd_0__inst_mult_12_180 ;
wire Xd_0__inst_mult_12_181 ;
wire Xd_0__inst_mult_12_182 ;
wire Xd_0__inst_mult_4_188 ;
wire Xd_0__inst_mult_4_189 ;
wire Xd_0__inst_mult_4_190 ;
wire Xd_0__inst_mult_9_173 ;
wire Xd_0__inst_mult_9_174 ;
wire Xd_0__inst_mult_9_175 ;
wire Xd_0__inst_mult_6_173 ;
wire Xd_0__inst_mult_6_174 ;
wire Xd_0__inst_mult_6_175 ;
wire Xd_0__inst_mult_14_188 ;
wire Xd_0__inst_mult_14_189 ;
wire Xd_0__inst_mult_14_190 ;
wire Xd_0__inst_mult_14_192 ;
wire Xd_0__inst_mult_14_193 ;
wire Xd_0__inst_mult_14_194 ;
wire Xd_0__inst_mult_8_177 ;
wire Xd_0__inst_mult_8_178 ;
wire Xd_0__inst_mult_8_179 ;
wire Xd_0__inst_mult_11_177 ;
wire Xd_0__inst_mult_11_178 ;
wire Xd_0__inst_mult_11_179 ;
wire Xd_0__inst_mult_10_173 ;
wire Xd_0__inst_mult_10_174 ;
wire Xd_0__inst_mult_10_175 ;
wire Xd_0__inst_mult_15_188 ;
wire Xd_0__inst_mult_15_189 ;
wire Xd_0__inst_mult_15_190 ;
wire Xd_0__inst_mult_13_177 ;
wire Xd_0__inst_mult_13_178 ;
wire Xd_0__inst_mult_13_179 ;
wire Xd_0__inst_mult_15_192 ;
wire Xd_0__inst_mult_15_193 ;
wire Xd_0__inst_mult_15_194 ;
wire Xd_0__inst_mult_12_184 ;
wire Xd_0__inst_mult_12_185 ;
wire Xd_0__inst_mult_12_186 ;
wire Xd_0__inst_mult_12_188 ;
wire Xd_0__inst_mult_12_189 ;
wire Xd_0__inst_mult_12_190 ;
wire Xd_0__inst_mult_4_192 ;
wire Xd_0__inst_mult_4_193 ;
wire Xd_0__inst_mult_4_194 ;
wire Xd_0__inst_mult_12_192 ;
wire Xd_0__inst_mult_12_193 ;
wire Xd_0__inst_mult_12_194 ;
wire Xd_0__inst_mult_13_180 ;
wire Xd_0__inst_mult_13_181 ;
wire Xd_0__inst_mult_13_182 ;
wire Xd_0__inst_mult_14_196 ;
wire Xd_0__inst_mult_14_197 ;
wire Xd_0__inst_mult_14_198 ;
wire Xd_0__inst_mult_15_196 ;
wire Xd_0__inst_mult_15_197 ;
wire Xd_0__inst_mult_15_198 ;
wire Xd_0__inst_mult_10_176 ;
wire Xd_0__inst_mult_10_177 ;
wire Xd_0__inst_mult_10_178 ;
wire Xd_0__inst_mult_11_180 ;
wire Xd_0__inst_mult_11_181 ;
wire Xd_0__inst_mult_11_182 ;
wire Xd_0__inst_mult_8_180 ;
wire Xd_0__inst_mult_8_181 ;
wire Xd_0__inst_mult_8_182 ;
wire Xd_0__inst_mult_9_176 ;
wire Xd_0__inst_mult_9_177 ;
wire Xd_0__inst_mult_9_178 ;
wire Xd_0__inst_mult_6_176 ;
wire Xd_0__inst_mult_6_177 ;
wire Xd_0__inst_mult_6_178 ;
wire Xd_0__inst_mult_7_169 ;
wire Xd_0__inst_mult_7_170 ;
wire Xd_0__inst_mult_7_171 ;
wire Xd_0__inst_mult_4_196 ;
wire Xd_0__inst_mult_4_197 ;
wire Xd_0__inst_mult_4_198 ;
wire Xd_0__inst_mult_5_169 ;
wire Xd_0__inst_mult_5_170 ;
wire Xd_0__inst_mult_5_171 ;
wire Xd_0__inst_mult_2_173 ;
wire Xd_0__inst_mult_2_174 ;
wire Xd_0__inst_mult_2_175 ;
wire Xd_0__inst_mult_3_169 ;
wire Xd_0__inst_mult_3_170 ;
wire Xd_0__inst_mult_3_171 ;
wire Xd_0__inst_mult_0_173 ;
wire Xd_0__inst_mult_0_174 ;
wire Xd_0__inst_mult_0_175 ;
wire Xd_0__inst_mult_1_173 ;
wire Xd_0__inst_mult_1_174 ;
wire Xd_0__inst_mult_1_175 ;
wire Xd_0__inst_mult_12_196 ;
wire Xd_0__inst_mult_12_197 ;
wire Xd_0__inst_mult_12_198 ;
wire Xd_0__inst_mult_13_184 ;
wire Xd_0__inst_mult_13_185 ;
wire Xd_0__inst_mult_13_186 ;
wire Xd_0__inst_mult_14_200 ;
wire Xd_0__inst_mult_14_201 ;
wire Xd_0__inst_mult_14_202 ;
wire Xd_0__inst_mult_15_200 ;
wire Xd_0__inst_mult_15_201 ;
wire Xd_0__inst_mult_15_202 ;
wire Xd_0__inst_mult_10_180 ;
wire Xd_0__inst_mult_10_181 ;
wire Xd_0__inst_mult_10_182 ;
wire Xd_0__inst_mult_11_184 ;
wire Xd_0__inst_mult_11_185 ;
wire Xd_0__inst_mult_11_186 ;
wire Xd_0__inst_mult_8_184 ;
wire Xd_0__inst_mult_8_185 ;
wire Xd_0__inst_mult_8_186 ;
wire Xd_0__inst_mult_9_180 ;
wire Xd_0__inst_mult_9_181 ;
wire Xd_0__inst_mult_9_182 ;
wire Xd_0__inst_mult_6_180 ;
wire Xd_0__inst_mult_6_181 ;
wire Xd_0__inst_mult_6_182 ;
wire Xd_0__inst_mult_7_173 ;
wire Xd_0__inst_mult_7_174 ;
wire Xd_0__inst_mult_7_175 ;
wire Xd_0__inst_mult_4_200 ;
wire Xd_0__inst_mult_4_201 ;
wire Xd_0__inst_mult_4_202 ;
wire Xd_0__inst_mult_5_173 ;
wire Xd_0__inst_mult_5_174 ;
wire Xd_0__inst_mult_5_175 ;
wire Xd_0__inst_mult_2_177 ;
wire Xd_0__inst_mult_2_178 ;
wire Xd_0__inst_mult_2_179 ;
wire Xd_0__inst_mult_3_173 ;
wire Xd_0__inst_mult_3_174 ;
wire Xd_0__inst_mult_3_175 ;
wire Xd_0__inst_mult_0_177 ;
wire Xd_0__inst_mult_0_178 ;
wire Xd_0__inst_mult_0_179 ;
wire Xd_0__inst_mult_1_177 ;
wire Xd_0__inst_mult_1_178 ;
wire Xd_0__inst_mult_1_179 ;
wire Xd_0__inst_mult_12_200 ;
wire Xd_0__inst_mult_12_201 ;
wire Xd_0__inst_mult_12_202 ;
wire Xd_0__inst_mult_13_188 ;
wire Xd_0__inst_mult_13_189 ;
wire Xd_0__inst_mult_13_190 ;
wire Xd_0__inst_mult_14_204 ;
wire Xd_0__inst_mult_14_205 ;
wire Xd_0__inst_mult_14_206 ;
wire Xd_0__inst_mult_15_204 ;
wire Xd_0__inst_mult_15_205 ;
wire Xd_0__inst_mult_15_206 ;
wire Xd_0__inst_mult_10_184 ;
wire Xd_0__inst_mult_10_185 ;
wire Xd_0__inst_mult_10_186 ;
wire Xd_0__inst_mult_11_188 ;
wire Xd_0__inst_mult_11_189 ;
wire Xd_0__inst_mult_11_190 ;
wire Xd_0__inst_mult_8_188 ;
wire Xd_0__inst_mult_8_189 ;
wire Xd_0__inst_mult_8_190 ;
wire Xd_0__inst_mult_9_184 ;
wire Xd_0__inst_mult_9_185 ;
wire Xd_0__inst_mult_9_186 ;
wire Xd_0__inst_mult_6_184 ;
wire Xd_0__inst_mult_6_185 ;
wire Xd_0__inst_mult_6_186 ;
wire Xd_0__inst_mult_7_176 ;
wire Xd_0__inst_mult_7_177 ;
wire Xd_0__inst_mult_7_178 ;
wire Xd_0__inst_mult_4_204 ;
wire Xd_0__inst_mult_4_205 ;
wire Xd_0__inst_mult_4_206 ;
wire Xd_0__inst_mult_5_176 ;
wire Xd_0__inst_mult_5_177 ;
wire Xd_0__inst_mult_5_178 ;
wire Xd_0__inst_mult_2_180 ;
wire Xd_0__inst_mult_2_181 ;
wire Xd_0__inst_mult_2_182 ;
wire Xd_0__inst_mult_3_176 ;
wire Xd_0__inst_mult_3_177 ;
wire Xd_0__inst_mult_3_178 ;
wire Xd_0__inst_mult_0_180 ;
wire Xd_0__inst_mult_0_181 ;
wire Xd_0__inst_mult_0_182 ;
wire Xd_0__inst_mult_1_180 ;
wire Xd_0__inst_mult_1_181 ;
wire Xd_0__inst_mult_1_182 ;
wire Xd_0__inst_mult_12_204 ;
wire Xd_0__inst_mult_12_205 ;
wire Xd_0__inst_mult_12_206 ;
wire Xd_0__inst_mult_13_192 ;
wire Xd_0__inst_mult_13_193 ;
wire Xd_0__inst_mult_13_194 ;
wire Xd_0__inst_mult_14_208 ;
wire Xd_0__inst_mult_14_209 ;
wire Xd_0__inst_mult_14_210 ;
wire Xd_0__inst_mult_15_208 ;
wire Xd_0__inst_mult_15_209 ;
wire Xd_0__inst_mult_15_210 ;
wire Xd_0__inst_mult_10_188 ;
wire Xd_0__inst_mult_10_189 ;
wire Xd_0__inst_mult_10_190 ;
wire Xd_0__inst_mult_11_192 ;
wire Xd_0__inst_mult_11_193 ;
wire Xd_0__inst_mult_11_194 ;
wire Xd_0__inst_mult_8_192 ;
wire Xd_0__inst_mult_8_193 ;
wire Xd_0__inst_mult_8_194 ;
wire Xd_0__inst_mult_9_188 ;
wire Xd_0__inst_mult_9_189 ;
wire Xd_0__inst_mult_9_190 ;
wire Xd_0__inst_mult_6_188 ;
wire Xd_0__inst_mult_6_189 ;
wire Xd_0__inst_mult_6_190 ;
wire Xd_0__inst_mult_7_180 ;
wire Xd_0__inst_mult_7_181 ;
wire Xd_0__inst_mult_7_182 ;
wire Xd_0__inst_mult_4_208 ;
wire Xd_0__inst_mult_4_209 ;
wire Xd_0__inst_mult_4_210 ;
wire Xd_0__inst_mult_5_180 ;
wire Xd_0__inst_mult_5_181 ;
wire Xd_0__inst_mult_5_182 ;
wire Xd_0__inst_mult_2_184 ;
wire Xd_0__inst_mult_2_185 ;
wire Xd_0__inst_mult_2_186 ;
wire Xd_0__inst_mult_3_180 ;
wire Xd_0__inst_mult_3_181 ;
wire Xd_0__inst_mult_3_182 ;
wire Xd_0__inst_mult_0_184 ;
wire Xd_0__inst_mult_0_185 ;
wire Xd_0__inst_mult_0_186 ;
wire Xd_0__inst_mult_1_184 ;
wire Xd_0__inst_mult_1_185 ;
wire Xd_0__inst_mult_1_186 ;
wire Xd_0__inst_mult_12_208 ;
wire Xd_0__inst_mult_12_209 ;
wire Xd_0__inst_mult_12_210 ;
wire Xd_0__inst_mult_13_196 ;
wire Xd_0__inst_mult_13_197 ;
wire Xd_0__inst_mult_13_198 ;
wire Xd_0__inst_mult_14_212 ;
wire Xd_0__inst_mult_14_213 ;
wire Xd_0__inst_mult_14_214 ;
wire Xd_0__inst_mult_15_212 ;
wire Xd_0__inst_mult_15_213 ;
wire Xd_0__inst_mult_15_214 ;
wire Xd_0__inst_mult_10_192 ;
wire Xd_0__inst_mult_10_193 ;
wire Xd_0__inst_mult_10_194 ;
wire Xd_0__inst_mult_11_196 ;
wire Xd_0__inst_mult_11_197 ;
wire Xd_0__inst_mult_11_198 ;
wire Xd_0__inst_mult_8_196 ;
wire Xd_0__inst_mult_8_197 ;
wire Xd_0__inst_mult_8_198 ;
wire Xd_0__inst_mult_9_192 ;
wire Xd_0__inst_mult_9_193 ;
wire Xd_0__inst_mult_9_194 ;
wire Xd_0__inst_mult_6_192 ;
wire Xd_0__inst_mult_6_193 ;
wire Xd_0__inst_mult_6_194 ;
wire Xd_0__inst_mult_7_184 ;
wire Xd_0__inst_mult_7_185 ;
wire Xd_0__inst_mult_7_186 ;
wire Xd_0__inst_mult_4_212 ;
wire Xd_0__inst_mult_4_213 ;
wire Xd_0__inst_mult_4_214 ;
wire Xd_0__inst_mult_5_184 ;
wire Xd_0__inst_mult_5_185 ;
wire Xd_0__inst_mult_5_186 ;
wire Xd_0__inst_mult_2_188 ;
wire Xd_0__inst_mult_2_189 ;
wire Xd_0__inst_mult_2_190 ;
wire Xd_0__inst_mult_3_184 ;
wire Xd_0__inst_mult_3_185 ;
wire Xd_0__inst_mult_3_186 ;
wire Xd_0__inst_mult_0_188 ;
wire Xd_0__inst_mult_0_189 ;
wire Xd_0__inst_mult_0_190 ;
wire Xd_0__inst_mult_1_188 ;
wire Xd_0__inst_mult_1_189 ;
wire Xd_0__inst_mult_1_190 ;
wire Xd_0__inst_mult_12_212 ;
wire Xd_0__inst_mult_12_213 ;
wire Xd_0__inst_mult_12_214 ;
wire Xd_0__inst_mult_13_200 ;
wire Xd_0__inst_mult_13_201 ;
wire Xd_0__inst_mult_13_202 ;
wire Xd_0__inst_mult_14_216 ;
wire Xd_0__inst_mult_14_217 ;
wire Xd_0__inst_mult_14_218 ;
wire Xd_0__inst_mult_15_216 ;
wire Xd_0__inst_mult_15_217 ;
wire Xd_0__inst_mult_15_218 ;
wire Xd_0__inst_mult_10_196 ;
wire Xd_0__inst_mult_10_197 ;
wire Xd_0__inst_mult_10_198 ;
wire Xd_0__inst_mult_11_200 ;
wire Xd_0__inst_mult_11_201 ;
wire Xd_0__inst_mult_11_202 ;
wire Xd_0__inst_mult_8_200 ;
wire Xd_0__inst_mult_8_201 ;
wire Xd_0__inst_mult_8_202 ;
wire Xd_0__inst_mult_9_196 ;
wire Xd_0__inst_mult_9_197 ;
wire Xd_0__inst_mult_9_198 ;
wire Xd_0__inst_mult_6_196 ;
wire Xd_0__inst_mult_6_197 ;
wire Xd_0__inst_mult_6_198 ;
wire Xd_0__inst_mult_7_188 ;
wire Xd_0__inst_mult_7_189 ;
wire Xd_0__inst_mult_7_190 ;
wire Xd_0__inst_mult_4_216 ;
wire Xd_0__inst_mult_4_217 ;
wire Xd_0__inst_mult_4_218 ;
wire Xd_0__inst_mult_5_188 ;
wire Xd_0__inst_mult_5_189 ;
wire Xd_0__inst_mult_5_190 ;
wire Xd_0__inst_mult_2_192 ;
wire Xd_0__inst_mult_2_193 ;
wire Xd_0__inst_mult_2_194 ;
wire Xd_0__inst_mult_3_188 ;
wire Xd_0__inst_mult_3_189 ;
wire Xd_0__inst_mult_3_190 ;
wire Xd_0__inst_mult_0_192 ;
wire Xd_0__inst_mult_0_193 ;
wire Xd_0__inst_mult_0_194 ;
wire Xd_0__inst_mult_1_192 ;
wire Xd_0__inst_mult_1_193 ;
wire Xd_0__inst_mult_1_194 ;
wire Xd_0__inst_mult_12_216 ;
wire Xd_0__inst_mult_12_217 ;
wire Xd_0__inst_mult_12_218 ;
wire Xd_0__inst_mult_13_204 ;
wire Xd_0__inst_mult_13_205 ;
wire Xd_0__inst_mult_13_206 ;
wire Xd_0__inst_mult_14_220 ;
wire Xd_0__inst_mult_14_221 ;
wire Xd_0__inst_mult_14_222 ;
wire Xd_0__inst_mult_15_220 ;
wire Xd_0__inst_mult_15_221 ;
wire Xd_0__inst_mult_15_222 ;
wire Xd_0__inst_mult_10_200 ;
wire Xd_0__inst_mult_10_201 ;
wire Xd_0__inst_mult_10_202 ;
wire Xd_0__inst_mult_11_204 ;
wire Xd_0__inst_mult_11_205 ;
wire Xd_0__inst_mult_11_206 ;
wire Xd_0__inst_mult_8_204 ;
wire Xd_0__inst_mult_8_205 ;
wire Xd_0__inst_mult_8_206 ;
wire Xd_0__inst_mult_9_200 ;
wire Xd_0__inst_mult_9_201 ;
wire Xd_0__inst_mult_9_202 ;
wire Xd_0__inst_mult_6_200 ;
wire Xd_0__inst_mult_6_201 ;
wire Xd_0__inst_mult_6_202 ;
wire Xd_0__inst_mult_7_192 ;
wire Xd_0__inst_mult_7_193 ;
wire Xd_0__inst_mult_7_194 ;
wire Xd_0__inst_mult_4_220 ;
wire Xd_0__inst_mult_4_221 ;
wire Xd_0__inst_mult_4_222 ;
wire Xd_0__inst_mult_5_192 ;
wire Xd_0__inst_mult_5_193 ;
wire Xd_0__inst_mult_5_194 ;
wire Xd_0__inst_mult_2_196 ;
wire Xd_0__inst_mult_2_197 ;
wire Xd_0__inst_mult_2_198 ;
wire Xd_0__inst_mult_3_192 ;
wire Xd_0__inst_mult_3_193 ;
wire Xd_0__inst_mult_3_194 ;
wire Xd_0__inst_mult_0_196 ;
wire Xd_0__inst_mult_0_197 ;
wire Xd_0__inst_mult_0_198 ;
wire Xd_0__inst_mult_1_196 ;
wire Xd_0__inst_mult_1_197 ;
wire Xd_0__inst_mult_1_198 ;
wire Xd_0__inst_mult_12_220 ;
wire Xd_0__inst_mult_12_221 ;
wire Xd_0__inst_mult_12_222 ;
wire Xd_0__inst_mult_13_208 ;
wire Xd_0__inst_mult_13_209 ;
wire Xd_0__inst_mult_13_210 ;
wire Xd_0__inst_mult_14_224 ;
wire Xd_0__inst_mult_14_225 ;
wire Xd_0__inst_mult_14_226 ;
wire Xd_0__inst_mult_15_224 ;
wire Xd_0__inst_mult_15_225 ;
wire Xd_0__inst_mult_15_226 ;
wire Xd_0__inst_mult_10_204 ;
wire Xd_0__inst_mult_10_205 ;
wire Xd_0__inst_mult_10_206 ;
wire Xd_0__inst_mult_11_208 ;
wire Xd_0__inst_mult_11_209 ;
wire Xd_0__inst_mult_11_210 ;
wire Xd_0__inst_mult_8_208 ;
wire Xd_0__inst_mult_8_209 ;
wire Xd_0__inst_mult_8_210 ;
wire Xd_0__inst_mult_9_204 ;
wire Xd_0__inst_mult_9_205 ;
wire Xd_0__inst_mult_9_206 ;
wire Xd_0__inst_mult_6_204 ;
wire Xd_0__inst_mult_6_205 ;
wire Xd_0__inst_mult_6_206 ;
wire Xd_0__inst_mult_7_196 ;
wire Xd_0__inst_mult_7_197 ;
wire Xd_0__inst_mult_7_198 ;
wire Xd_0__inst_mult_4_224 ;
wire Xd_0__inst_mult_4_225 ;
wire Xd_0__inst_mult_4_226 ;
wire Xd_0__inst_mult_5_196 ;
wire Xd_0__inst_mult_5_197 ;
wire Xd_0__inst_mult_5_198 ;
wire Xd_0__inst_mult_2_200 ;
wire Xd_0__inst_mult_2_201 ;
wire Xd_0__inst_mult_2_202 ;
wire Xd_0__inst_mult_3_196 ;
wire Xd_0__inst_mult_3_197 ;
wire Xd_0__inst_mult_3_198 ;
wire Xd_0__inst_mult_0_200 ;
wire Xd_0__inst_mult_0_201 ;
wire Xd_0__inst_mult_0_202 ;
wire Xd_0__inst_mult_1_200 ;
wire Xd_0__inst_mult_1_201 ;
wire Xd_0__inst_mult_1_202 ;
wire Xd_0__inst_mult_12_224 ;
wire Xd_0__inst_mult_12_225 ;
wire Xd_0__inst_mult_12_226 ;
wire Xd_0__inst_mult_13_212 ;
wire Xd_0__inst_mult_13_213 ;
wire Xd_0__inst_mult_13_214 ;
wire Xd_0__inst_mult_14_228 ;
wire Xd_0__inst_mult_14_229 ;
wire Xd_0__inst_mult_14_230 ;
wire Xd_0__inst_mult_15_228 ;
wire Xd_0__inst_mult_15_229 ;
wire Xd_0__inst_mult_15_230 ;
wire Xd_0__inst_mult_10_208 ;
wire Xd_0__inst_mult_10_209 ;
wire Xd_0__inst_mult_10_210 ;
wire Xd_0__inst_mult_11_212 ;
wire Xd_0__inst_mult_11_213 ;
wire Xd_0__inst_mult_11_214 ;
wire Xd_0__inst_mult_8_212 ;
wire Xd_0__inst_mult_8_213 ;
wire Xd_0__inst_mult_8_214 ;
wire Xd_0__inst_mult_9_208 ;
wire Xd_0__inst_mult_9_209 ;
wire Xd_0__inst_mult_9_210 ;
wire Xd_0__inst_mult_6_208 ;
wire Xd_0__inst_mult_6_209 ;
wire Xd_0__inst_mult_6_210 ;
wire Xd_0__inst_mult_7_200 ;
wire Xd_0__inst_mult_7_201 ;
wire Xd_0__inst_mult_7_202 ;
wire Xd_0__inst_mult_4_228 ;
wire Xd_0__inst_mult_4_229 ;
wire Xd_0__inst_mult_4_230 ;
wire Xd_0__inst_mult_5_200 ;
wire Xd_0__inst_mult_5_201 ;
wire Xd_0__inst_mult_5_202 ;
wire Xd_0__inst_mult_2_204 ;
wire Xd_0__inst_mult_2_205 ;
wire Xd_0__inst_mult_2_206 ;
wire Xd_0__inst_mult_3_200 ;
wire Xd_0__inst_mult_3_201 ;
wire Xd_0__inst_mult_3_202 ;
wire Xd_0__inst_mult_0_204 ;
wire Xd_0__inst_mult_0_205 ;
wire Xd_0__inst_mult_0_206 ;
wire Xd_0__inst_mult_1_204 ;
wire Xd_0__inst_mult_1_205 ;
wire Xd_0__inst_mult_1_206 ;
wire Xd_0__inst_mult_12_228 ;
wire Xd_0__inst_mult_12_229 ;
wire Xd_0__inst_mult_12_230 ;
wire Xd_0__inst_mult_13_216 ;
wire Xd_0__inst_mult_13_217 ;
wire Xd_0__inst_mult_13_218 ;
wire Xd_0__inst_mult_14_232 ;
wire Xd_0__inst_mult_14_233 ;
wire Xd_0__inst_mult_14_234 ;
wire Xd_0__inst_mult_15_232 ;
wire Xd_0__inst_mult_15_233 ;
wire Xd_0__inst_mult_15_234 ;
wire Xd_0__inst_mult_10_212 ;
wire Xd_0__inst_mult_10_213 ;
wire Xd_0__inst_mult_10_214 ;
wire Xd_0__inst_mult_11_216 ;
wire Xd_0__inst_mult_11_217 ;
wire Xd_0__inst_mult_11_218 ;
wire Xd_0__inst_mult_8_216 ;
wire Xd_0__inst_mult_8_217 ;
wire Xd_0__inst_mult_8_218 ;
wire Xd_0__inst_mult_9_212 ;
wire Xd_0__inst_mult_9_213 ;
wire Xd_0__inst_mult_9_214 ;
wire Xd_0__inst_mult_6_212 ;
wire Xd_0__inst_mult_6_213 ;
wire Xd_0__inst_mult_6_214 ;
wire Xd_0__inst_mult_7_204 ;
wire Xd_0__inst_mult_7_205 ;
wire Xd_0__inst_mult_7_206 ;
wire Xd_0__inst_mult_4_232 ;
wire Xd_0__inst_mult_4_233 ;
wire Xd_0__inst_mult_4_234 ;
wire Xd_0__inst_mult_5_204 ;
wire Xd_0__inst_mult_5_205 ;
wire Xd_0__inst_mult_5_206 ;
wire Xd_0__inst_mult_2_208 ;
wire Xd_0__inst_mult_2_209 ;
wire Xd_0__inst_mult_2_210 ;
wire Xd_0__inst_mult_3_204 ;
wire Xd_0__inst_mult_3_205 ;
wire Xd_0__inst_mult_3_206 ;
wire Xd_0__inst_mult_0_208 ;
wire Xd_0__inst_mult_0_209 ;
wire Xd_0__inst_mult_0_210 ;
wire Xd_0__inst_mult_1_208 ;
wire Xd_0__inst_mult_1_209 ;
wire Xd_0__inst_mult_1_210 ;
wire Xd_0__inst_mult_12_232 ;
wire Xd_0__inst_mult_12_233 ;
wire Xd_0__inst_mult_12_234 ;
wire Xd_0__inst_mult_13_220 ;
wire Xd_0__inst_mult_13_221 ;
wire Xd_0__inst_mult_13_222 ;
wire Xd_0__inst_mult_14_236 ;
wire Xd_0__inst_mult_14_237 ;
wire Xd_0__inst_mult_14_238 ;
wire Xd_0__inst_mult_15_236 ;
wire Xd_0__inst_mult_15_237 ;
wire Xd_0__inst_mult_15_238 ;
wire Xd_0__inst_mult_10_216 ;
wire Xd_0__inst_mult_10_217 ;
wire Xd_0__inst_mult_10_218 ;
wire Xd_0__inst_mult_11_220 ;
wire Xd_0__inst_mult_11_221 ;
wire Xd_0__inst_mult_11_222 ;
wire Xd_0__inst_mult_8_220 ;
wire Xd_0__inst_mult_8_221 ;
wire Xd_0__inst_mult_8_222 ;
wire Xd_0__inst_mult_9_216 ;
wire Xd_0__inst_mult_9_217 ;
wire Xd_0__inst_mult_9_218 ;
wire Xd_0__inst_mult_6_216 ;
wire Xd_0__inst_mult_6_217 ;
wire Xd_0__inst_mult_6_218 ;
wire Xd_0__inst_mult_7_208 ;
wire Xd_0__inst_mult_7_209 ;
wire Xd_0__inst_mult_7_210 ;
wire Xd_0__inst_mult_4_236 ;
wire Xd_0__inst_mult_4_237 ;
wire Xd_0__inst_mult_4_238 ;
wire Xd_0__inst_mult_5_208 ;
wire Xd_0__inst_mult_5_209 ;
wire Xd_0__inst_mult_5_210 ;
wire Xd_0__inst_mult_2_212 ;
wire Xd_0__inst_mult_2_213 ;
wire Xd_0__inst_mult_2_214 ;
wire Xd_0__inst_mult_3_208 ;
wire Xd_0__inst_mult_3_209 ;
wire Xd_0__inst_mult_3_210 ;
wire Xd_0__inst_mult_0_212 ;
wire Xd_0__inst_mult_0_213 ;
wire Xd_0__inst_mult_0_214 ;
wire Xd_0__inst_mult_1_212 ;
wire Xd_0__inst_mult_1_213 ;
wire Xd_0__inst_mult_1_214 ;
wire Xd_0__inst_mult_12_236 ;
wire Xd_0__inst_mult_12_237 ;
wire Xd_0__inst_mult_12_238 ;
wire Xd_0__inst_mult_13_224 ;
wire Xd_0__inst_mult_13_225 ;
wire Xd_0__inst_mult_13_226 ;
wire Xd_0__inst_mult_14_240 ;
wire Xd_0__inst_mult_14_241 ;
wire Xd_0__inst_mult_14_242 ;
wire Xd_0__inst_mult_15_240 ;
wire Xd_0__inst_mult_15_241 ;
wire Xd_0__inst_mult_15_242 ;
wire Xd_0__inst_mult_10_220 ;
wire Xd_0__inst_mult_10_221 ;
wire Xd_0__inst_mult_10_222 ;
wire Xd_0__inst_mult_11_224 ;
wire Xd_0__inst_mult_11_225 ;
wire Xd_0__inst_mult_11_226 ;
wire Xd_0__inst_mult_8_224 ;
wire Xd_0__inst_mult_8_225 ;
wire Xd_0__inst_mult_8_226 ;
wire Xd_0__inst_mult_9_220 ;
wire Xd_0__inst_mult_9_221 ;
wire Xd_0__inst_mult_9_222 ;
wire Xd_0__inst_mult_6_220 ;
wire Xd_0__inst_mult_6_221 ;
wire Xd_0__inst_mult_6_222 ;
wire Xd_0__inst_mult_7_212 ;
wire Xd_0__inst_mult_7_213 ;
wire Xd_0__inst_mult_7_214 ;
wire Xd_0__inst_mult_4_240 ;
wire Xd_0__inst_mult_4_241 ;
wire Xd_0__inst_mult_4_242 ;
wire Xd_0__inst_mult_5_212 ;
wire Xd_0__inst_mult_5_213 ;
wire Xd_0__inst_mult_5_214 ;
wire Xd_0__inst_mult_2_216 ;
wire Xd_0__inst_mult_2_217 ;
wire Xd_0__inst_mult_2_218 ;
wire Xd_0__inst_mult_3_212 ;
wire Xd_0__inst_mult_3_213 ;
wire Xd_0__inst_mult_3_214 ;
wire Xd_0__inst_mult_0_216 ;
wire Xd_0__inst_mult_0_217 ;
wire Xd_0__inst_mult_0_218 ;
wire Xd_0__inst_mult_1_216 ;
wire Xd_0__inst_mult_1_217 ;
wire Xd_0__inst_mult_1_218 ;
wire Xd_0__inst_mult_12_240 ;
wire Xd_0__inst_mult_12_241 ;
wire Xd_0__inst_mult_12_242 ;
wire Xd_0__inst_mult_13_228 ;
wire Xd_0__inst_mult_13_229 ;
wire Xd_0__inst_mult_13_230 ;
wire Xd_0__inst_mult_14_244 ;
wire Xd_0__inst_mult_14_245 ;
wire Xd_0__inst_mult_14_246 ;
wire Xd_0__inst_mult_15_244 ;
wire Xd_0__inst_mult_15_245 ;
wire Xd_0__inst_mult_15_246 ;
wire Xd_0__inst_mult_10_224 ;
wire Xd_0__inst_mult_10_225 ;
wire Xd_0__inst_mult_10_226 ;
wire Xd_0__inst_mult_11_228 ;
wire Xd_0__inst_mult_11_229 ;
wire Xd_0__inst_mult_11_230 ;
wire Xd_0__inst_mult_8_228 ;
wire Xd_0__inst_mult_8_229 ;
wire Xd_0__inst_mult_8_230 ;
wire Xd_0__inst_mult_9_224 ;
wire Xd_0__inst_mult_9_225 ;
wire Xd_0__inst_mult_9_226 ;
wire Xd_0__inst_mult_6_224 ;
wire Xd_0__inst_mult_6_225 ;
wire Xd_0__inst_mult_6_226 ;
wire Xd_0__inst_mult_7_216 ;
wire Xd_0__inst_mult_7_217 ;
wire Xd_0__inst_mult_7_218 ;
wire Xd_0__inst_mult_4_244 ;
wire Xd_0__inst_mult_4_245 ;
wire Xd_0__inst_mult_4_246 ;
wire Xd_0__inst_mult_5_216 ;
wire Xd_0__inst_mult_5_217 ;
wire Xd_0__inst_mult_5_218 ;
wire Xd_0__inst_mult_2_220 ;
wire Xd_0__inst_mult_2_221 ;
wire Xd_0__inst_mult_2_222 ;
wire Xd_0__inst_mult_3_216 ;
wire Xd_0__inst_mult_3_217 ;
wire Xd_0__inst_mult_3_218 ;
wire Xd_0__inst_mult_0_220 ;
wire Xd_0__inst_mult_0_221 ;
wire Xd_0__inst_mult_0_222 ;
wire Xd_0__inst_mult_1_220 ;
wire Xd_0__inst_mult_1_221 ;
wire Xd_0__inst_mult_1_222 ;
wire Xd_0__inst_mult_12_244 ;
wire Xd_0__inst_mult_12_245 ;
wire Xd_0__inst_mult_12_246 ;
wire Xd_0__inst_mult_13_232 ;
wire Xd_0__inst_mult_13_233 ;
wire Xd_0__inst_mult_13_234 ;
wire Xd_0__inst_mult_14_248 ;
wire Xd_0__inst_mult_14_249 ;
wire Xd_0__inst_mult_14_250 ;
wire Xd_0__inst_mult_15_248 ;
wire Xd_0__inst_mult_15_249 ;
wire Xd_0__inst_mult_15_250 ;
wire Xd_0__inst_mult_10_228 ;
wire Xd_0__inst_mult_10_229 ;
wire Xd_0__inst_mult_10_230 ;
wire Xd_0__inst_mult_11_232 ;
wire Xd_0__inst_mult_11_233 ;
wire Xd_0__inst_mult_11_234 ;
wire Xd_0__inst_mult_8_232 ;
wire Xd_0__inst_mult_8_233 ;
wire Xd_0__inst_mult_8_234 ;
wire Xd_0__inst_mult_9_228 ;
wire Xd_0__inst_mult_9_229 ;
wire Xd_0__inst_mult_9_230 ;
wire Xd_0__inst_mult_6_228 ;
wire Xd_0__inst_mult_6_229 ;
wire Xd_0__inst_mult_6_230 ;
wire Xd_0__inst_mult_7_220 ;
wire Xd_0__inst_mult_7_221 ;
wire Xd_0__inst_mult_7_222 ;
wire Xd_0__inst_mult_4_248 ;
wire Xd_0__inst_mult_4_249 ;
wire Xd_0__inst_mult_4_250 ;
wire Xd_0__inst_mult_5_220 ;
wire Xd_0__inst_mult_5_221 ;
wire Xd_0__inst_mult_5_222 ;
wire Xd_0__inst_mult_2_224 ;
wire Xd_0__inst_mult_2_225 ;
wire Xd_0__inst_mult_2_226 ;
wire Xd_0__inst_mult_3_220 ;
wire Xd_0__inst_mult_3_221 ;
wire Xd_0__inst_mult_3_222 ;
wire Xd_0__inst_mult_0_224 ;
wire Xd_0__inst_mult_0_225 ;
wire Xd_0__inst_mult_0_226 ;
wire Xd_0__inst_mult_1_224 ;
wire Xd_0__inst_mult_1_225 ;
wire Xd_0__inst_mult_1_226 ;
wire Xd_0__inst_mult_12_248 ;
wire Xd_0__inst_mult_12_249 ;
wire Xd_0__inst_mult_12_250 ;
wire Xd_0__inst_mult_13_236 ;
wire Xd_0__inst_mult_13_237 ;
wire Xd_0__inst_mult_13_238 ;
wire Xd_0__inst_mult_14_252 ;
wire Xd_0__inst_mult_14_253 ;
wire Xd_0__inst_mult_14_254 ;
wire Xd_0__inst_mult_15_252 ;
wire Xd_0__inst_mult_15_253 ;
wire Xd_0__inst_mult_15_254 ;
wire Xd_0__inst_mult_10_232 ;
wire Xd_0__inst_mult_10_233 ;
wire Xd_0__inst_mult_10_234 ;
wire Xd_0__inst_mult_11_236 ;
wire Xd_0__inst_mult_11_237 ;
wire Xd_0__inst_mult_11_238 ;
wire Xd_0__inst_mult_8_236 ;
wire Xd_0__inst_mult_8_237 ;
wire Xd_0__inst_mult_8_238 ;
wire Xd_0__inst_mult_9_232 ;
wire Xd_0__inst_mult_9_233 ;
wire Xd_0__inst_mult_9_234 ;
wire Xd_0__inst_mult_6_232 ;
wire Xd_0__inst_mult_6_233 ;
wire Xd_0__inst_mult_6_234 ;
wire Xd_0__inst_mult_7_224 ;
wire Xd_0__inst_mult_7_225 ;
wire Xd_0__inst_mult_7_226 ;
wire Xd_0__inst_mult_4_252 ;
wire Xd_0__inst_mult_4_253 ;
wire Xd_0__inst_mult_4_254 ;
wire Xd_0__inst_mult_5_224 ;
wire Xd_0__inst_mult_5_225 ;
wire Xd_0__inst_mult_5_226 ;
wire Xd_0__inst_mult_2_228 ;
wire Xd_0__inst_mult_2_229 ;
wire Xd_0__inst_mult_2_230 ;
wire Xd_0__inst_mult_3_224 ;
wire Xd_0__inst_mult_3_225 ;
wire Xd_0__inst_mult_3_226 ;
wire Xd_0__inst_mult_0_228 ;
wire Xd_0__inst_mult_0_229 ;
wire Xd_0__inst_mult_0_230 ;
wire Xd_0__inst_mult_1_228 ;
wire Xd_0__inst_mult_1_229 ;
wire Xd_0__inst_mult_1_230 ;
wire Xd_0__inst_mult_12_252 ;
wire Xd_0__inst_mult_12_253 ;
wire Xd_0__inst_mult_12_254 ;
wire Xd_0__inst_mult_13_240 ;
wire Xd_0__inst_mult_13_241 ;
wire Xd_0__inst_mult_13_242 ;
wire Xd_0__inst_mult_14_256 ;
wire Xd_0__inst_mult_14_257 ;
wire Xd_0__inst_mult_14_258 ;
wire Xd_0__inst_mult_15_256 ;
wire Xd_0__inst_mult_15_257 ;
wire Xd_0__inst_mult_15_258 ;
wire Xd_0__inst_mult_10_236 ;
wire Xd_0__inst_mult_10_237 ;
wire Xd_0__inst_mult_10_238 ;
wire Xd_0__inst_mult_11_240 ;
wire Xd_0__inst_mult_11_241 ;
wire Xd_0__inst_mult_11_242 ;
wire Xd_0__inst_mult_8_240 ;
wire Xd_0__inst_mult_8_241 ;
wire Xd_0__inst_mult_8_242 ;
wire Xd_0__inst_mult_9_236 ;
wire Xd_0__inst_mult_9_237 ;
wire Xd_0__inst_mult_9_238 ;
wire Xd_0__inst_mult_6_236 ;
wire Xd_0__inst_mult_6_237 ;
wire Xd_0__inst_mult_6_238 ;
wire Xd_0__inst_mult_7_228 ;
wire Xd_0__inst_mult_7_229 ;
wire Xd_0__inst_mult_7_230 ;
wire Xd_0__inst_mult_4_256 ;
wire Xd_0__inst_mult_4_257 ;
wire Xd_0__inst_mult_4_258 ;
wire Xd_0__inst_mult_5_228 ;
wire Xd_0__inst_mult_5_229 ;
wire Xd_0__inst_mult_5_230 ;
wire Xd_0__inst_mult_2_232 ;
wire Xd_0__inst_mult_2_233 ;
wire Xd_0__inst_mult_2_234 ;
wire Xd_0__inst_mult_3_228 ;
wire Xd_0__inst_mult_3_229 ;
wire Xd_0__inst_mult_3_230 ;
wire Xd_0__inst_mult_0_232 ;
wire Xd_0__inst_mult_0_233 ;
wire Xd_0__inst_mult_0_234 ;
wire Xd_0__inst_mult_1_232 ;
wire Xd_0__inst_mult_1_233 ;
wire Xd_0__inst_mult_1_234 ;
wire Xd_0__inst_mult_12_256 ;
wire Xd_0__inst_mult_13_244 ;
wire Xd_0__inst_mult_14_260 ;
wire Xd_0__inst_mult_15_260 ;
wire Xd_0__inst_mult_10_240 ;
wire Xd_0__inst_mult_11_244 ;
wire Xd_0__inst_mult_8_244 ;
wire Xd_0__inst_mult_9_240 ;
wire Xd_0__inst_mult_6_240 ;
wire Xd_0__inst_mult_7_232 ;
wire Xd_0__inst_mult_4_260 ;
wire Xd_0__inst_mult_5_232 ;
wire Xd_0__inst_mult_2_236 ;
wire Xd_0__inst_mult_3_232 ;
wire Xd_0__inst_mult_0_236 ;
wire Xd_0__inst_mult_1_236 ;
wire Xd_0__inst_mult_12_260 ;
wire Xd_0__inst_mult_12_261 ;
wire Xd_0__inst_mult_12_262 ;
wire Xd_0__inst_mult_13_248 ;
wire Xd_0__inst_mult_13_249 ;
wire Xd_0__inst_mult_13_250 ;
wire Xd_0__inst_i29_1_sumout ;
wire Xd_0__inst_i29_2 ;
wire Xd_0__inst_i29_3 ;
wire Xd_0__inst_i29_5_sumout ;
wire Xd_0__inst_i29_6 ;
wire Xd_0__inst_i29_7 ;
wire Xd_0__inst_mult_9_244 ;
wire Xd_0__inst_mult_9_248 ;
wire Xd_0__inst_mult_9_249 ;
wire Xd_0__inst_mult_9_250 ;
wire Xd_0__inst_mult_14_264 ;
wire Xd_0__inst_mult_14_265 ;
wire Xd_0__inst_mult_14_266 ;
wire Xd_0__inst_mult_15_264 ;
wire Xd_0__inst_mult_15_265 ;
wire Xd_0__inst_mult_15_266 ;
wire Xd_0__inst_i29_9_sumout ;
wire Xd_0__inst_i29_10 ;
wire Xd_0__inst_i29_11 ;
wire Xd_0__inst_i29_13_sumout ;
wire Xd_0__inst_i29_14 ;
wire Xd_0__inst_i29_15 ;
wire Xd_0__inst_mult_6_244 ;
wire Xd_0__inst_mult_6_248 ;
wire Xd_0__inst_mult_6_249 ;
wire Xd_0__inst_mult_6_250 ;
wire Xd_0__inst_mult_14_268 ;
wire Xd_0__inst_mult_14_269 ;
wire Xd_0__inst_mult_14_270 ;
wire Xd_0__inst_mult_14_272 ;
wire Xd_0__inst_mult_14_276 ;
wire Xd_0__inst_mult_14_277 ;
wire Xd_0__inst_mult_14_278 ;
wire Xd_0__inst_mult_10_244 ;
wire Xd_0__inst_mult_10_245 ;
wire Xd_0__inst_mult_10_246 ;
wire Xd_0__inst_mult_11_248 ;
wire Xd_0__inst_mult_11_249 ;
wire Xd_0__inst_mult_11_250 ;
wire Xd_0__inst_i29_17_sumout ;
wire Xd_0__inst_i29_18 ;
wire Xd_0__inst_i29_19 ;
wire Xd_0__inst_i29_21_sumout ;
wire Xd_0__inst_i29_22 ;
wire Xd_0__inst_i29_23 ;
wire Xd_0__inst_mult_8_248 ;
wire Xd_0__inst_mult_8_252 ;
wire Xd_0__inst_mult_8_253 ;
wire Xd_0__inst_mult_8_254 ;
wire Xd_0__inst_mult_8_256 ;
wire Xd_0__inst_mult_8_257 ;
wire Xd_0__inst_mult_8_258 ;
wire Xd_0__inst_mult_9_252 ;
wire Xd_0__inst_mult_9_253 ;
wire Xd_0__inst_mult_9_254 ;
wire Xd_0__inst_i29_25_sumout ;
wire Xd_0__inst_i29_26 ;
wire Xd_0__inst_i29_27 ;
wire Xd_0__inst_i29_29_sumout ;
wire Xd_0__inst_i29_30 ;
wire Xd_0__inst_i29_31 ;
wire Xd_0__inst_mult_11_252 ;
wire Xd_0__inst_mult_11_256 ;
wire Xd_0__inst_mult_11_257 ;
wire Xd_0__inst_mult_11_258 ;
wire Xd_0__inst_mult_6_252 ;
wire Xd_0__inst_mult_6_253 ;
wire Xd_0__inst_mult_6_254 ;
wire Xd_0__inst_mult_7_236 ;
wire Xd_0__inst_mult_7_237 ;
wire Xd_0__inst_mult_7_238 ;
wire Xd_0__inst_i29_33_sumout ;
wire Xd_0__inst_i29_34 ;
wire Xd_0__inst_i29_35 ;
wire Xd_0__inst_i29_37_sumout ;
wire Xd_0__inst_i29_38 ;
wire Xd_0__inst_i29_39 ;
wire Xd_0__inst_mult_10_248 ;
wire Xd_0__inst_mult_10_252 ;
wire Xd_0__inst_mult_10_253 ;
wire Xd_0__inst_mult_10_254 ;
wire Xd_0__inst_mult_15_268 ;
wire Xd_0__inst_mult_15_269 ;
wire Xd_0__inst_mult_15_270 ;
wire Xd_0__inst_mult_4_264 ;
wire Xd_0__inst_mult_4_265 ;
wire Xd_0__inst_mult_4_266 ;
wire Xd_0__inst_mult_5_236 ;
wire Xd_0__inst_mult_5_237 ;
wire Xd_0__inst_mult_5_238 ;
wire Xd_0__inst_i29_41_sumout ;
wire Xd_0__inst_i29_42 ;
wire Xd_0__inst_i29_43 ;
wire Xd_0__inst_i29_45_sumout ;
wire Xd_0__inst_i29_46 ;
wire Xd_0__inst_i29_47 ;
wire Xd_0__inst_mult_13_252 ;
wire Xd_0__inst_mult_13_256 ;
wire Xd_0__inst_mult_13_257 ;
wire Xd_0__inst_mult_13_258 ;
wire Xd_0__inst_mult_2_240 ;
wire Xd_0__inst_mult_2_241 ;
wire Xd_0__inst_mult_2_242 ;
wire Xd_0__inst_mult_3_236 ;
wire Xd_0__inst_mult_3_237 ;
wire Xd_0__inst_mult_3_238 ;
wire Xd_0__inst_i29_49_sumout ;
wire Xd_0__inst_i29_50 ;
wire Xd_0__inst_i29_51 ;
wire Xd_0__inst_i29_53_sumout ;
wire Xd_0__inst_i29_54 ;
wire Xd_0__inst_i29_55 ;
wire Xd_0__inst_mult_15_272 ;
wire Xd_0__inst_mult_15_276 ;
wire Xd_0__inst_mult_15_277 ;
wire Xd_0__inst_mult_15_278 ;
wire Xd_0__inst_mult_0_240 ;
wire Xd_0__inst_mult_0_241 ;
wire Xd_0__inst_mult_0_242 ;
wire Xd_0__inst_mult_1_240 ;
wire Xd_0__inst_mult_1_241 ;
wire Xd_0__inst_mult_1_242 ;
wire Xd_0__inst_i29_57_sumout ;
wire Xd_0__inst_i29_58 ;
wire Xd_0__inst_i29_59 ;
wire Xd_0__inst_i29_61_sumout ;
wire Xd_0__inst_i29_62 ;
wire Xd_0__inst_i29_63 ;
wire Xd_0__inst_mult_12_264 ;
wire Xd_0__inst_mult_12_268 ;
wire Xd_0__inst_mult_12_269 ;
wire Xd_0__inst_mult_12_270 ;
wire Xd_0__inst_mult_12_272 ;
wire Xd_0__inst_mult_12_273 ;
wire Xd_0__inst_mult_12_274 ;
wire Xd_0__inst_mult_4_268 ;
wire Xd_0__inst_mult_4_269 ;
wire Xd_0__inst_mult_4_270 ;
wire Xd_0__inst_mult_12_276 ;
wire Xd_0__inst_mult_12_277 ;
wire Xd_0__inst_mult_12_278 ;
wire Xd_0__inst_mult_13_260 ;
wire Xd_0__inst_mult_13_261 ;
wire Xd_0__inst_mult_13_262 ;
wire Xd_0__inst_mult_14_280 ;
wire Xd_0__inst_mult_14_281 ;
wire Xd_0__inst_mult_14_282 ;
wire Xd_0__inst_mult_15_280 ;
wire Xd_0__inst_mult_15_281 ;
wire Xd_0__inst_mult_15_282 ;
wire Xd_0__inst_mult_10_256 ;
wire Xd_0__inst_mult_10_257 ;
wire Xd_0__inst_mult_10_258 ;
wire Xd_0__inst_mult_11_260 ;
wire Xd_0__inst_mult_11_261 ;
wire Xd_0__inst_mult_11_262 ;
wire Xd_0__inst_mult_8_260 ;
wire Xd_0__inst_mult_8_261 ;
wire Xd_0__inst_mult_8_262 ;
wire Xd_0__inst_mult_9_256 ;
wire Xd_0__inst_mult_9_257 ;
wire Xd_0__inst_mult_9_258 ;
wire Xd_0__inst_mult_6_256 ;
wire Xd_0__inst_mult_6_257 ;
wire Xd_0__inst_mult_6_258 ;
wire Xd_0__inst_mult_7_240 ;
wire Xd_0__inst_mult_7_241 ;
wire Xd_0__inst_mult_7_242 ;
wire Xd_0__inst_mult_4_272 ;
wire Xd_0__inst_mult_4_273 ;
wire Xd_0__inst_mult_4_274 ;
wire Xd_0__inst_mult_5_240 ;
wire Xd_0__inst_mult_5_241 ;
wire Xd_0__inst_mult_5_242 ;
wire Xd_0__inst_mult_2_244 ;
wire Xd_0__inst_mult_2_245 ;
wire Xd_0__inst_mult_2_246 ;
wire Xd_0__inst_mult_3_240 ;
wire Xd_0__inst_mult_3_241 ;
wire Xd_0__inst_mult_3_242 ;
wire Xd_0__inst_mult_0_244 ;
wire Xd_0__inst_mult_0_245 ;
wire Xd_0__inst_mult_0_246 ;
wire Xd_0__inst_mult_1_244 ;
wire Xd_0__inst_mult_1_245 ;
wire Xd_0__inst_mult_1_246 ;
wire Xd_0__inst_mult_12_280 ;
wire Xd_0__inst_mult_12_281 ;
wire Xd_0__inst_mult_12_282 ;
wire Xd_0__inst_mult_13_264 ;
wire Xd_0__inst_mult_13_265 ;
wire Xd_0__inst_mult_13_266 ;
wire Xd_0__inst_mult_14_284 ;
wire Xd_0__inst_mult_14_285 ;
wire Xd_0__inst_mult_14_286 ;
wire Xd_0__inst_mult_15_284 ;
wire Xd_0__inst_mult_15_285 ;
wire Xd_0__inst_mult_15_286 ;
wire Xd_0__inst_mult_10_260 ;
wire Xd_0__inst_mult_10_261 ;
wire Xd_0__inst_mult_10_262 ;
wire Xd_0__inst_mult_11_264 ;
wire Xd_0__inst_mult_11_265 ;
wire Xd_0__inst_mult_11_266 ;
wire Xd_0__inst_mult_8_264 ;
wire Xd_0__inst_mult_8_265 ;
wire Xd_0__inst_mult_8_266 ;
wire Xd_0__inst_mult_9_260 ;
wire Xd_0__inst_mult_9_261 ;
wire Xd_0__inst_mult_9_262 ;
wire Xd_0__inst_mult_6_260 ;
wire Xd_0__inst_mult_6_261 ;
wire Xd_0__inst_mult_6_262 ;
wire Xd_0__inst_mult_7_244 ;
wire Xd_0__inst_mult_7_245 ;
wire Xd_0__inst_mult_7_246 ;
wire Xd_0__inst_mult_4_276 ;
wire Xd_0__inst_mult_4_277 ;
wire Xd_0__inst_mult_4_278 ;
wire Xd_0__inst_mult_5_244 ;
wire Xd_0__inst_mult_5_245 ;
wire Xd_0__inst_mult_5_246 ;
wire Xd_0__inst_mult_2_248 ;
wire Xd_0__inst_mult_2_249 ;
wire Xd_0__inst_mult_2_250 ;
wire Xd_0__inst_mult_3_244 ;
wire Xd_0__inst_mult_3_245 ;
wire Xd_0__inst_mult_3_246 ;
wire Xd_0__inst_mult_0_248 ;
wire Xd_0__inst_mult_0_249 ;
wire Xd_0__inst_mult_0_250 ;
wire Xd_0__inst_mult_1_248 ;
wire Xd_0__inst_mult_1_249 ;
wire Xd_0__inst_mult_1_250 ;
wire Xd_0__inst_mult_12_284 ;
wire Xd_0__inst_mult_12_285 ;
wire Xd_0__inst_mult_12_286 ;
wire Xd_0__inst_mult_13_268 ;
wire Xd_0__inst_mult_13_269 ;
wire Xd_0__inst_mult_13_270 ;
wire Xd_0__inst_mult_14_288 ;
wire Xd_0__inst_mult_14_289 ;
wire Xd_0__inst_mult_14_290 ;
wire Xd_0__inst_mult_15_288 ;
wire Xd_0__inst_mult_15_289 ;
wire Xd_0__inst_mult_15_290 ;
wire Xd_0__inst_mult_10_264 ;
wire Xd_0__inst_mult_10_265 ;
wire Xd_0__inst_mult_10_266 ;
wire Xd_0__inst_mult_11_268 ;
wire Xd_0__inst_mult_11_269 ;
wire Xd_0__inst_mult_11_270 ;
wire Xd_0__inst_mult_8_268 ;
wire Xd_0__inst_mult_8_269 ;
wire Xd_0__inst_mult_8_270 ;
wire Xd_0__inst_mult_9_264 ;
wire Xd_0__inst_mult_9_265 ;
wire Xd_0__inst_mult_9_266 ;
wire Xd_0__inst_mult_6_264 ;
wire Xd_0__inst_mult_6_265 ;
wire Xd_0__inst_mult_6_266 ;
wire Xd_0__inst_mult_7_248 ;
wire Xd_0__inst_mult_7_249 ;
wire Xd_0__inst_mult_7_250 ;
wire Xd_0__inst_mult_4_280 ;
wire Xd_0__inst_mult_4_281 ;
wire Xd_0__inst_mult_4_282 ;
wire Xd_0__inst_mult_5_248 ;
wire Xd_0__inst_mult_5_249 ;
wire Xd_0__inst_mult_5_250 ;
wire Xd_0__inst_mult_2_252 ;
wire Xd_0__inst_mult_2_253 ;
wire Xd_0__inst_mult_2_254 ;
wire Xd_0__inst_mult_3_248 ;
wire Xd_0__inst_mult_3_249 ;
wire Xd_0__inst_mult_3_250 ;
wire Xd_0__inst_mult_0_252 ;
wire Xd_0__inst_mult_0_253 ;
wire Xd_0__inst_mult_0_254 ;
wire Xd_0__inst_mult_1_252 ;
wire Xd_0__inst_mult_1_253 ;
wire Xd_0__inst_mult_1_254 ;
wire Xd_0__inst_mult_12_288 ;
wire Xd_0__inst_mult_12_289 ;
wire Xd_0__inst_mult_12_290 ;
wire Xd_0__inst_mult_13_272 ;
wire Xd_0__inst_mult_13_273 ;
wire Xd_0__inst_mult_13_274 ;
wire Xd_0__inst_mult_14_292 ;
wire Xd_0__inst_mult_14_293 ;
wire Xd_0__inst_mult_14_294 ;
wire Xd_0__inst_mult_15_292 ;
wire Xd_0__inst_mult_15_293 ;
wire Xd_0__inst_mult_15_294 ;
wire Xd_0__inst_mult_10_268 ;
wire Xd_0__inst_mult_10_269 ;
wire Xd_0__inst_mult_10_270 ;
wire Xd_0__inst_mult_11_272 ;
wire Xd_0__inst_mult_11_273 ;
wire Xd_0__inst_mult_11_274 ;
wire Xd_0__inst_mult_8_272 ;
wire Xd_0__inst_mult_8_273 ;
wire Xd_0__inst_mult_8_274 ;
wire Xd_0__inst_mult_9_268 ;
wire Xd_0__inst_mult_9_269 ;
wire Xd_0__inst_mult_9_270 ;
wire Xd_0__inst_mult_6_268 ;
wire Xd_0__inst_mult_6_269 ;
wire Xd_0__inst_mult_6_270 ;
wire Xd_0__inst_mult_7_252 ;
wire Xd_0__inst_mult_7_253 ;
wire Xd_0__inst_mult_7_254 ;
wire Xd_0__inst_mult_4_284 ;
wire Xd_0__inst_mult_4_285 ;
wire Xd_0__inst_mult_4_286 ;
wire Xd_0__inst_mult_5_252 ;
wire Xd_0__inst_mult_5_253 ;
wire Xd_0__inst_mult_5_254 ;
wire Xd_0__inst_mult_2_256 ;
wire Xd_0__inst_mult_2_257 ;
wire Xd_0__inst_mult_2_258 ;
wire Xd_0__inst_mult_3_252 ;
wire Xd_0__inst_mult_3_253 ;
wire Xd_0__inst_mult_3_254 ;
wire Xd_0__inst_mult_0_256 ;
wire Xd_0__inst_mult_0_257 ;
wire Xd_0__inst_mult_0_258 ;
wire Xd_0__inst_mult_1_256 ;
wire Xd_0__inst_mult_1_257 ;
wire Xd_0__inst_mult_1_258 ;
wire Xd_0__inst_mult_12_35_sumout ;
wire Xd_0__inst_mult_12_36 ;
wire Xd_0__inst_mult_12_37 ;
wire Xd_0__inst_mult_1_35_sumout ;
wire Xd_0__inst_mult_1_36 ;
wire Xd_0__inst_mult_1_37 ;
wire Xd_0__inst_mult_6_35_sumout ;
wire Xd_0__inst_mult_6_36 ;
wire Xd_0__inst_mult_6_37 ;
wire Xd_0__inst_mult_5_35_sumout ;
wire Xd_0__inst_mult_5_36 ;
wire Xd_0__inst_mult_5_37 ;
wire Xd_0__inst_mult_2_35_sumout ;
wire Xd_0__inst_mult_2_36 ;
wire Xd_0__inst_mult_2_37 ;
wire Xd_0__inst_mult_14_35_sumout ;
wire Xd_0__inst_mult_14_36 ;
wire Xd_0__inst_mult_14_37 ;
wire Xd_0__inst_mult_12_39_sumout ;
wire Xd_0__inst_mult_12_40 ;
wire Xd_0__inst_mult_12_41 ;
wire Xd_0__inst_mult_15_35_sumout ;
wire Xd_0__inst_mult_15_36 ;
wire Xd_0__inst_mult_15_37 ;
wire Xd_0__inst_mult_5_39_sumout ;
wire Xd_0__inst_mult_5_40 ;
wire Xd_0__inst_mult_5_41 ;
wire Xd_0__inst_mult_4_35_sumout ;
wire Xd_0__inst_mult_4_36 ;
wire Xd_0__inst_mult_4_37 ;
wire Xd_0__inst_mult_10_35_sumout ;
wire Xd_0__inst_mult_10_36 ;
wire Xd_0__inst_mult_10_37 ;
wire Xd_0__inst_mult_6_39_sumout ;
wire Xd_0__inst_mult_6_40 ;
wire Xd_0__inst_mult_6_41 ;
wire Xd_0__inst_mult_2_39_sumout ;
wire Xd_0__inst_mult_2_40 ;
wire Xd_0__inst_mult_2_41 ;
wire Xd_0__inst_mult_13_35_sumout ;
wire Xd_0__inst_mult_13_36 ;
wire Xd_0__inst_mult_13_37 ;
wire Xd_0__inst_mult_14_39_sumout ;
wire Xd_0__inst_mult_14_40 ;
wire Xd_0__inst_mult_14_41 ;
wire Xd_0__inst_mult_3_35_sumout ;
wire Xd_0__inst_mult_3_36 ;
wire Xd_0__inst_mult_3_37 ;
wire Xd_0__inst_mult_9_272 ;
wire Xd_0__inst_mult_9_273 ;
wire Xd_0__inst_mult_9_274 ;
wire Xd_0__inst_mult_9_276 ;
wire Xd_0__inst_mult_9_277 ;
wire Xd_0__inst_mult_9_278 ;
wire Xd_0__inst_mult_14_43_sumout ;
wire Xd_0__inst_mult_14_44 ;
wire Xd_0__inst_mult_14_45 ;
wire Xd_0__inst_mult_6_272 ;
wire Xd_0__inst_mult_6_273 ;
wire Xd_0__inst_mult_6_274 ;
wire Xd_0__inst_mult_6_276 ;
wire Xd_0__inst_mult_6_277 ;
wire Xd_0__inst_mult_6_278 ;
wire Xd_0__inst_mult_14_296 ;
wire Xd_0__inst_mult_14_297 ;
wire Xd_0__inst_mult_14_298 ;
wire Xd_0__inst_mult_14_300 ;
wire Xd_0__inst_mult_14_301 ;
wire Xd_0__inst_mult_14_302 ;
wire Xd_0__inst_mult_14_304 ;
wire Xd_0__inst_mult_14_305 ;
wire Xd_0__inst_mult_14_306 ;
wire Xd_0__inst_mult_8_276 ;
wire Xd_0__inst_mult_8_277 ;
wire Xd_0__inst_mult_8_278 ;
wire Xd_0__inst_mult_8_280 ;
wire Xd_0__inst_mult_8_281 ;
wire Xd_0__inst_mult_8_282 ;
wire Xd_0__inst_mult_9_35_sumout ;
wire Xd_0__inst_mult_9_36 ;
wire Xd_0__inst_mult_9_37 ;
wire Xd_0__inst_mult_11_276 ;
wire Xd_0__inst_mult_11_277 ;
wire Xd_0__inst_mult_11_278 ;
wire Xd_0__inst_mult_11_280 ;
wire Xd_0__inst_mult_11_281 ;
wire Xd_0__inst_mult_11_282 ;
wire Xd_0__inst_mult_10_272 ;
wire Xd_0__inst_mult_10_273 ;
wire Xd_0__inst_mult_10_274 ;
wire Xd_0__inst_mult_10_276 ;
wire Xd_0__inst_mult_10_277 ;
wire Xd_0__inst_mult_10_278 ;
wire Xd_0__inst_mult_15_296 ;
wire Xd_0__inst_mult_15_297 ;
wire Xd_0__inst_mult_15_298 ;
wire Xd_0__inst_mult_13_276 ;
wire Xd_0__inst_mult_13_277 ;
wire Xd_0__inst_mult_13_278 ;
wire Xd_0__inst_mult_13_280 ;
wire Xd_0__inst_mult_13_281 ;
wire Xd_0__inst_mult_13_282 ;
wire Xd_0__inst_mult_15_300 ;
wire Xd_0__inst_mult_15_301 ;
wire Xd_0__inst_mult_15_302 ;
wire Xd_0__inst_mult_15_304 ;
wire Xd_0__inst_mult_15_305 ;
wire Xd_0__inst_mult_15_306 ;
wire Xd_0__inst_mult_12_292 ;
wire Xd_0__inst_mult_12_293 ;
wire Xd_0__inst_mult_12_294 ;
wire Xd_0__inst_mult_12_296 ;
wire Xd_0__inst_mult_12_297 ;
wire Xd_0__inst_mult_12_298 ;
wire Xd_0__inst_mult_12_300 ;
wire Xd_0__inst_mult_12_301 ;
wire Xd_0__inst_mult_12_302 ;
wire Xd_0__inst_mult_4_288 ;
wire Xd_0__inst_mult_4_289 ;
wire Xd_0__inst_mult_4_290 ;
wire Xd_0__inst_mult_12_305 ;
wire Xd_0__inst_mult_12_306 ;
wire Xd_0__inst_mult_13_285 ;
wire Xd_0__inst_mult_13_286 ;
wire Xd_0__inst_mult_14_309 ;
wire Xd_0__inst_mult_14_310 ;
wire Xd_0__inst_mult_15_309 ;
wire Xd_0__inst_mult_15_310 ;
wire Xd_0__inst_mult_10_281 ;
wire Xd_0__inst_mult_10_282 ;
wire Xd_0__inst_mult_11_285 ;
wire Xd_0__inst_mult_11_286 ;
wire Xd_0__inst_mult_8_285 ;
wire Xd_0__inst_mult_8_286 ;
wire Xd_0__inst_mult_9_281 ;
wire Xd_0__inst_mult_9_282 ;
wire Xd_0__inst_mult_6_281 ;
wire Xd_0__inst_mult_6_282 ;
wire Xd_0__inst_mult_7_257 ;
wire Xd_0__inst_mult_7_258 ;
wire Xd_0__inst_mult_4_293 ;
wire Xd_0__inst_mult_4_294 ;
wire Xd_0__inst_mult_5_257 ;
wire Xd_0__inst_mult_5_258 ;
wire Xd_0__inst_mult_2_261 ;
wire Xd_0__inst_mult_2_262 ;
wire Xd_0__inst_mult_3_257 ;
wire Xd_0__inst_mult_3_258 ;
wire Xd_0__inst_mult_0_261 ;
wire Xd_0__inst_mult_0_262 ;
wire Xd_0__inst_mult_1_261 ;
wire Xd_0__inst_mult_1_262 ;
wire Xd_0__inst_mult_12_308 ;
wire Xd_0__inst_mult_12_309 ;
wire Xd_0__inst_mult_12_310 ;
wire Xd_0__inst_mult_12_312 ;
wire Xd_0__inst_mult_12_313 ;
wire Xd_0__inst_mult_12_314 ;
wire Xd_0__inst_mult_13_288 ;
wire Xd_0__inst_mult_13_289 ;
wire Xd_0__inst_mult_13_290 ;
wire Xd_0__inst_mult_13_292 ;
wire Xd_0__inst_mult_13_293 ;
wire Xd_0__inst_mult_13_294 ;
wire Xd_0__inst_mult_14_312 ;
wire Xd_0__inst_mult_14_313 ;
wire Xd_0__inst_mult_14_314 ;
wire Xd_0__inst_mult_14_316 ;
wire Xd_0__inst_mult_14_317 ;
wire Xd_0__inst_mult_14_318 ;
wire Xd_0__inst_mult_15_312 ;
wire Xd_0__inst_mult_15_313 ;
wire Xd_0__inst_mult_15_314 ;
wire Xd_0__inst_mult_15_316 ;
wire Xd_0__inst_mult_15_317 ;
wire Xd_0__inst_mult_15_318 ;
wire Xd_0__inst_mult_10_284 ;
wire Xd_0__inst_mult_10_285 ;
wire Xd_0__inst_mult_10_286 ;
wire Xd_0__inst_mult_10_288 ;
wire Xd_0__inst_mult_10_289 ;
wire Xd_0__inst_mult_10_290 ;
wire Xd_0__inst_mult_11_288 ;
wire Xd_0__inst_mult_11_289 ;
wire Xd_0__inst_mult_11_290 ;
wire Xd_0__inst_mult_11_292 ;
wire Xd_0__inst_mult_11_293 ;
wire Xd_0__inst_mult_11_294 ;
wire Xd_0__inst_mult_8_288 ;
wire Xd_0__inst_mult_8_289 ;
wire Xd_0__inst_mult_8_290 ;
wire Xd_0__inst_mult_8_292 ;
wire Xd_0__inst_mult_8_293 ;
wire Xd_0__inst_mult_8_294 ;
wire Xd_0__inst_mult_9_284 ;
wire Xd_0__inst_mult_9_285 ;
wire Xd_0__inst_mult_9_286 ;
wire Xd_0__inst_mult_9_288 ;
wire Xd_0__inst_mult_9_289 ;
wire Xd_0__inst_mult_9_290 ;
wire Xd_0__inst_mult_6_284 ;
wire Xd_0__inst_mult_6_285 ;
wire Xd_0__inst_mult_6_286 ;
wire Xd_0__inst_mult_6_288 ;
wire Xd_0__inst_mult_6_289 ;
wire Xd_0__inst_mult_6_290 ;
wire Xd_0__inst_mult_7_260 ;
wire Xd_0__inst_mult_7_261 ;
wire Xd_0__inst_mult_7_262 ;
wire Xd_0__inst_mult_7_264 ;
wire Xd_0__inst_mult_7_265 ;
wire Xd_0__inst_mult_7_266 ;
wire Xd_0__inst_mult_4_296 ;
wire Xd_0__inst_mult_4_297 ;
wire Xd_0__inst_mult_4_298 ;
wire Xd_0__inst_mult_4_300 ;
wire Xd_0__inst_mult_4_301 ;
wire Xd_0__inst_mult_4_302 ;
wire Xd_0__inst_mult_5_260 ;
wire Xd_0__inst_mult_5_261 ;
wire Xd_0__inst_mult_5_262 ;
wire Xd_0__inst_mult_5_264 ;
wire Xd_0__inst_mult_5_265 ;
wire Xd_0__inst_mult_5_266 ;
wire Xd_0__inst_mult_2_264 ;
wire Xd_0__inst_mult_2_265 ;
wire Xd_0__inst_mult_2_266 ;
wire Xd_0__inst_mult_2_268 ;
wire Xd_0__inst_mult_2_269 ;
wire Xd_0__inst_mult_2_270 ;
wire Xd_0__inst_mult_3_260 ;
wire Xd_0__inst_mult_3_261 ;
wire Xd_0__inst_mult_3_262 ;
wire Xd_0__inst_mult_3_264 ;
wire Xd_0__inst_mult_3_265 ;
wire Xd_0__inst_mult_3_266 ;
wire Xd_0__inst_mult_0_264 ;
wire Xd_0__inst_mult_0_265 ;
wire Xd_0__inst_mult_0_266 ;
wire Xd_0__inst_mult_0_268 ;
wire Xd_0__inst_mult_0_269 ;
wire Xd_0__inst_mult_0_270 ;
wire Xd_0__inst_mult_1_264 ;
wire Xd_0__inst_mult_1_265 ;
wire Xd_0__inst_mult_1_266 ;
wire Xd_0__inst_mult_1_268 ;
wire Xd_0__inst_mult_1_269 ;
wire Xd_0__inst_mult_1_270 ;
wire Xd_0__inst_mult_12_316 ;
wire Xd_0__inst_mult_12_317 ;
wire Xd_0__inst_mult_12_318 ;
wire Xd_0__inst_mult_12_320 ;
wire Xd_0__inst_mult_12_321 ;
wire Xd_0__inst_mult_12_322 ;
wire Xd_0__inst_mult_13_39_sumout ;
wire Xd_0__inst_mult_13_40 ;
wire Xd_0__inst_mult_13_41 ;
wire Xd_0__inst_mult_13_296 ;
wire Xd_0__inst_mult_13_297 ;
wire Xd_0__inst_mult_13_298 ;
wire Xd_0__inst_mult_13_300 ;
wire Xd_0__inst_mult_13_301 ;
wire Xd_0__inst_mult_13_302 ;
wire Xd_0__inst_mult_14_47_sumout ;
wire Xd_0__inst_mult_14_48 ;
wire Xd_0__inst_mult_14_49 ;
wire Xd_0__inst_mult_14_320 ;
wire Xd_0__inst_mult_14_321 ;
wire Xd_0__inst_mult_14_322 ;
wire Xd_0__inst_mult_14_324 ;
wire Xd_0__inst_mult_14_325 ;
wire Xd_0__inst_mult_14_326 ;
wire Xd_0__inst_mult_7_35_sumout ;
wire Xd_0__inst_mult_7_36 ;
wire Xd_0__inst_mult_7_37 ;
wire Xd_0__inst_mult_15_320 ;
wire Xd_0__inst_mult_15_321 ;
wire Xd_0__inst_mult_15_322 ;
wire Xd_0__inst_mult_15_324 ;
wire Xd_0__inst_mult_15_325 ;
wire Xd_0__inst_mult_15_326 ;
wire Xd_0__inst_mult_8_35_sumout ;
wire Xd_0__inst_mult_8_36 ;
wire Xd_0__inst_mult_8_37 ;
wire Xd_0__inst_mult_10_292 ;
wire Xd_0__inst_mult_10_293 ;
wire Xd_0__inst_mult_10_294 ;
wire Xd_0__inst_mult_10_296 ;
wire Xd_0__inst_mult_10_297 ;
wire Xd_0__inst_mult_10_298 ;
wire Xd_0__inst_mult_3_39_sumout ;
wire Xd_0__inst_mult_3_40 ;
wire Xd_0__inst_mult_3_41 ;
wire Xd_0__inst_mult_11_296 ;
wire Xd_0__inst_mult_11_297 ;
wire Xd_0__inst_mult_11_298 ;
wire Xd_0__inst_mult_11_300 ;
wire Xd_0__inst_mult_11_301 ;
wire Xd_0__inst_mult_11_302 ;
wire Xd_0__inst_mult_15_39_sumout ;
wire Xd_0__inst_mult_15_40 ;
wire Xd_0__inst_mult_15_41 ;
wire Xd_0__inst_mult_8_296 ;
wire Xd_0__inst_mult_8_297 ;
wire Xd_0__inst_mult_8_298 ;
wire Xd_0__inst_mult_8_300 ;
wire Xd_0__inst_mult_8_301 ;
wire Xd_0__inst_mult_8_302 ;
wire Xd_0__inst_mult_3_43_sumout ;
wire Xd_0__inst_mult_3_44 ;
wire Xd_0__inst_mult_3_45 ;
wire Xd_0__inst_mult_9_292 ;
wire Xd_0__inst_mult_9_293 ;
wire Xd_0__inst_mult_9_294 ;
wire Xd_0__inst_mult_9_296 ;
wire Xd_0__inst_mult_9_297 ;
wire Xd_0__inst_mult_9_298 ;
wire Xd_0__inst_mult_1_39_sumout ;
wire Xd_0__inst_mult_1_40 ;
wire Xd_0__inst_mult_1_41 ;
wire Xd_0__inst_mult_6_292 ;
wire Xd_0__inst_mult_6_293 ;
wire Xd_0__inst_mult_6_294 ;
wire Xd_0__inst_mult_6_296 ;
wire Xd_0__inst_mult_6_297 ;
wire Xd_0__inst_mult_6_298 ;
wire Xd_0__inst_mult_12_43_sumout ;
wire Xd_0__inst_mult_12_44 ;
wire Xd_0__inst_mult_12_45 ;
wire Xd_0__inst_mult_7_268 ;
wire Xd_0__inst_mult_7_269 ;
wire Xd_0__inst_mult_7_270 ;
wire Xd_0__inst_mult_7_272 ;
wire Xd_0__inst_mult_7_273 ;
wire Xd_0__inst_mult_7_274 ;
wire Xd_0__inst_mult_11_35_sumout ;
wire Xd_0__inst_mult_11_36 ;
wire Xd_0__inst_mult_11_37 ;
wire Xd_0__inst_mult_4_304 ;
wire Xd_0__inst_mult_4_305 ;
wire Xd_0__inst_mult_4_306 ;
wire Xd_0__inst_mult_4_308 ;
wire Xd_0__inst_mult_4_309 ;
wire Xd_0__inst_mult_4_310 ;
wire Xd_0__inst_mult_8_39_sumout ;
wire Xd_0__inst_mult_8_40 ;
wire Xd_0__inst_mult_8_41 ;
wire Xd_0__inst_mult_5_268 ;
wire Xd_0__inst_mult_5_269 ;
wire Xd_0__inst_mult_5_270 ;
wire Xd_0__inst_mult_5_272 ;
wire Xd_0__inst_mult_5_273 ;
wire Xd_0__inst_mult_5_274 ;
wire Xd_0__inst_mult_8_43_sumout ;
wire Xd_0__inst_mult_8_44 ;
wire Xd_0__inst_mult_8_45 ;
wire Xd_0__inst_mult_2_272 ;
wire Xd_0__inst_mult_2_273 ;
wire Xd_0__inst_mult_2_274 ;
wire Xd_0__inst_mult_2_276 ;
wire Xd_0__inst_mult_2_277 ;
wire Xd_0__inst_mult_2_278 ;
wire Xd_0__inst_mult_14_51_sumout ;
wire Xd_0__inst_mult_14_52 ;
wire Xd_0__inst_mult_14_53 ;
wire Xd_0__inst_mult_3_268 ;
wire Xd_0__inst_mult_3_269 ;
wire Xd_0__inst_mult_3_270 ;
wire Xd_0__inst_mult_3_272 ;
wire Xd_0__inst_mult_3_273 ;
wire Xd_0__inst_mult_3_274 ;
wire Xd_0__inst_mult_10_39_sumout ;
wire Xd_0__inst_mult_10_40 ;
wire Xd_0__inst_mult_10_41 ;
wire Xd_0__inst_mult_0_272 ;
wire Xd_0__inst_mult_0_273 ;
wire Xd_0__inst_mult_0_274 ;
wire Xd_0__inst_mult_0_276 ;
wire Xd_0__inst_mult_0_277 ;
wire Xd_0__inst_mult_0_278 ;
wire Xd_0__inst_mult_15_43_sumout ;
wire Xd_0__inst_mult_15_44 ;
wire Xd_0__inst_mult_15_45 ;
wire Xd_0__inst_mult_1_272 ;
wire Xd_0__inst_mult_1_273 ;
wire Xd_0__inst_mult_1_274 ;
wire Xd_0__inst_mult_1_276 ;
wire Xd_0__inst_mult_1_277 ;
wire Xd_0__inst_mult_1_278 ;
wire Xd_0__inst_mult_0_35_sumout ;
wire Xd_0__inst_mult_0_36 ;
wire Xd_0__inst_mult_0_37 ;
wire Xd_0__inst_mult_12_324 ;
wire Xd_0__inst_mult_12_325 ;
wire Xd_0__inst_mult_12_326 ;
wire Xd_0__inst_mult_12_328 ;
wire Xd_0__inst_mult_12_329 ;
wire Xd_0__inst_mult_12_330 ;
wire Xd_0__inst_mult_13_304 ;
wire Xd_0__inst_mult_13_305 ;
wire Xd_0__inst_mult_13_306 ;
wire Xd_0__inst_mult_13_308 ;
wire Xd_0__inst_mult_13_309 ;
wire Xd_0__inst_mult_13_310 ;
wire Xd_0__inst_mult_14_328 ;
wire Xd_0__inst_mult_14_329 ;
wire Xd_0__inst_mult_14_330 ;
wire Xd_0__inst_mult_14_332 ;
wire Xd_0__inst_mult_14_333 ;
wire Xd_0__inst_mult_14_334 ;
wire Xd_0__inst_mult_15_328 ;
wire Xd_0__inst_mult_15_329 ;
wire Xd_0__inst_mult_15_330 ;
wire Xd_0__inst_mult_15_332 ;
wire Xd_0__inst_mult_15_333 ;
wire Xd_0__inst_mult_15_334 ;
wire Xd_0__inst_mult_10_300 ;
wire Xd_0__inst_mult_10_301 ;
wire Xd_0__inst_mult_10_302 ;
wire Xd_0__inst_mult_10_304 ;
wire Xd_0__inst_mult_10_305 ;
wire Xd_0__inst_mult_10_306 ;
wire Xd_0__inst_mult_11_304 ;
wire Xd_0__inst_mult_11_305 ;
wire Xd_0__inst_mult_11_306 ;
wire Xd_0__inst_mult_11_308 ;
wire Xd_0__inst_mult_11_309 ;
wire Xd_0__inst_mult_11_310 ;
wire Xd_0__inst_mult_8_304 ;
wire Xd_0__inst_mult_8_305 ;
wire Xd_0__inst_mult_8_306 ;
wire Xd_0__inst_mult_8_308 ;
wire Xd_0__inst_mult_8_309 ;
wire Xd_0__inst_mult_8_310 ;
wire Xd_0__inst_mult_9_300 ;
wire Xd_0__inst_mult_9_301 ;
wire Xd_0__inst_mult_9_302 ;
wire Xd_0__inst_mult_9_304 ;
wire Xd_0__inst_mult_9_305 ;
wire Xd_0__inst_mult_9_306 ;
wire Xd_0__inst_mult_6_300 ;
wire Xd_0__inst_mult_6_301 ;
wire Xd_0__inst_mult_6_302 ;
wire Xd_0__inst_mult_6_304 ;
wire Xd_0__inst_mult_6_305 ;
wire Xd_0__inst_mult_6_306 ;
wire Xd_0__inst_mult_7_276 ;
wire Xd_0__inst_mult_7_277 ;
wire Xd_0__inst_mult_7_278 ;
wire Xd_0__inst_mult_7_280 ;
wire Xd_0__inst_mult_7_281 ;
wire Xd_0__inst_mult_7_282 ;
wire Xd_0__inst_mult_4_312 ;
wire Xd_0__inst_mult_4_313 ;
wire Xd_0__inst_mult_4_314 ;
wire Xd_0__inst_mult_4_316 ;
wire Xd_0__inst_mult_4_317 ;
wire Xd_0__inst_mult_4_318 ;
wire Xd_0__inst_mult_5_276 ;
wire Xd_0__inst_mult_5_277 ;
wire Xd_0__inst_mult_5_278 ;
wire Xd_0__inst_mult_5_280 ;
wire Xd_0__inst_mult_5_281 ;
wire Xd_0__inst_mult_5_282 ;
wire Xd_0__inst_mult_2_280 ;
wire Xd_0__inst_mult_2_281 ;
wire Xd_0__inst_mult_2_282 ;
wire Xd_0__inst_mult_2_284 ;
wire Xd_0__inst_mult_2_285 ;
wire Xd_0__inst_mult_2_286 ;
wire Xd_0__inst_mult_3_276 ;
wire Xd_0__inst_mult_3_277 ;
wire Xd_0__inst_mult_3_278 ;
wire Xd_0__inst_mult_3_280 ;
wire Xd_0__inst_mult_3_281 ;
wire Xd_0__inst_mult_3_282 ;
wire Xd_0__inst_mult_0_280 ;
wire Xd_0__inst_mult_0_281 ;
wire Xd_0__inst_mult_0_282 ;
wire Xd_0__inst_mult_0_284 ;
wire Xd_0__inst_mult_0_285 ;
wire Xd_0__inst_mult_0_286 ;
wire Xd_0__inst_mult_1_280 ;
wire Xd_0__inst_mult_1_281 ;
wire Xd_0__inst_mult_1_282 ;
wire Xd_0__inst_mult_1_284 ;
wire Xd_0__inst_mult_1_285 ;
wire Xd_0__inst_mult_1_286 ;
wire Xd_0__inst_mult_12_332 ;
wire Xd_0__inst_mult_12_333 ;
wire Xd_0__inst_mult_12_334 ;
wire Xd_0__inst_mult_12_336 ;
wire Xd_0__inst_mult_12_337 ;
wire Xd_0__inst_mult_12_338 ;
wire Xd_0__inst_mult_13_312 ;
wire Xd_0__inst_mult_13_313 ;
wire Xd_0__inst_mult_13_314 ;
wire Xd_0__inst_mult_13_316 ;
wire Xd_0__inst_mult_13_317 ;
wire Xd_0__inst_mult_13_318 ;
wire Xd_0__inst_mult_14_336 ;
wire Xd_0__inst_mult_14_337 ;
wire Xd_0__inst_mult_14_338 ;
wire Xd_0__inst_mult_14_340 ;
wire Xd_0__inst_mult_14_341 ;
wire Xd_0__inst_mult_14_342 ;
wire Xd_0__inst_mult_15_336 ;
wire Xd_0__inst_mult_15_337 ;
wire Xd_0__inst_mult_15_338 ;
wire Xd_0__inst_mult_15_340 ;
wire Xd_0__inst_mult_15_341 ;
wire Xd_0__inst_mult_15_342 ;
wire Xd_0__inst_mult_10_308 ;
wire Xd_0__inst_mult_10_309 ;
wire Xd_0__inst_mult_10_310 ;
wire Xd_0__inst_mult_10_312 ;
wire Xd_0__inst_mult_10_313 ;
wire Xd_0__inst_mult_10_314 ;
wire Xd_0__inst_mult_11_312 ;
wire Xd_0__inst_mult_11_313 ;
wire Xd_0__inst_mult_11_314 ;
wire Xd_0__inst_mult_11_316 ;
wire Xd_0__inst_mult_11_317 ;
wire Xd_0__inst_mult_11_318 ;
wire Xd_0__inst_mult_8_312 ;
wire Xd_0__inst_mult_8_313 ;
wire Xd_0__inst_mult_8_314 ;
wire Xd_0__inst_mult_8_316 ;
wire Xd_0__inst_mult_8_317 ;
wire Xd_0__inst_mult_8_318 ;
wire Xd_0__inst_mult_9_308 ;
wire Xd_0__inst_mult_9_309 ;
wire Xd_0__inst_mult_9_310 ;
wire Xd_0__inst_mult_9_312 ;
wire Xd_0__inst_mult_9_313 ;
wire Xd_0__inst_mult_9_314 ;
wire Xd_0__inst_mult_6_308 ;
wire Xd_0__inst_mult_6_309 ;
wire Xd_0__inst_mult_6_310 ;
wire Xd_0__inst_mult_6_312 ;
wire Xd_0__inst_mult_6_313 ;
wire Xd_0__inst_mult_6_314 ;
wire Xd_0__inst_mult_7_284 ;
wire Xd_0__inst_mult_7_285 ;
wire Xd_0__inst_mult_7_286 ;
wire Xd_0__inst_mult_7_288 ;
wire Xd_0__inst_mult_7_289 ;
wire Xd_0__inst_mult_7_290 ;
wire Xd_0__inst_mult_4_320 ;
wire Xd_0__inst_mult_4_321 ;
wire Xd_0__inst_mult_4_322 ;
wire Xd_0__inst_mult_4_324 ;
wire Xd_0__inst_mult_4_325 ;
wire Xd_0__inst_mult_4_326 ;
wire Xd_0__inst_mult_5_284 ;
wire Xd_0__inst_mult_5_285 ;
wire Xd_0__inst_mult_5_286 ;
wire Xd_0__inst_mult_5_288 ;
wire Xd_0__inst_mult_5_289 ;
wire Xd_0__inst_mult_5_290 ;
wire Xd_0__inst_mult_2_288 ;
wire Xd_0__inst_mult_2_289 ;
wire Xd_0__inst_mult_2_290 ;
wire Xd_0__inst_mult_2_292 ;
wire Xd_0__inst_mult_2_293 ;
wire Xd_0__inst_mult_2_294 ;
wire Xd_0__inst_mult_3_284 ;
wire Xd_0__inst_mult_3_285 ;
wire Xd_0__inst_mult_3_286 ;
wire Xd_0__inst_mult_3_288 ;
wire Xd_0__inst_mult_3_289 ;
wire Xd_0__inst_mult_3_290 ;
wire Xd_0__inst_mult_0_288 ;
wire Xd_0__inst_mult_0_289 ;
wire Xd_0__inst_mult_0_290 ;
wire Xd_0__inst_mult_0_292 ;
wire Xd_0__inst_mult_0_293 ;
wire Xd_0__inst_mult_0_294 ;
wire Xd_0__inst_mult_1_288 ;
wire Xd_0__inst_mult_1_289 ;
wire Xd_0__inst_mult_1_290 ;
wire Xd_0__inst_mult_1_292 ;
wire Xd_0__inst_mult_1_293 ;
wire Xd_0__inst_mult_1_294 ;
wire Xd_0__inst_mult_12_340 ;
wire Xd_0__inst_mult_12_341 ;
wire Xd_0__inst_mult_12_342 ;
wire Xd_0__inst_mult_12_344 ;
wire Xd_0__inst_mult_12_345 ;
wire Xd_0__inst_mult_12_346 ;
wire Xd_0__inst_mult_13_320 ;
wire Xd_0__inst_mult_13_321 ;
wire Xd_0__inst_mult_13_322 ;
wire Xd_0__inst_mult_13_324 ;
wire Xd_0__inst_mult_13_325 ;
wire Xd_0__inst_mult_13_326 ;
wire Xd_0__inst_mult_14_344 ;
wire Xd_0__inst_mult_14_345 ;
wire Xd_0__inst_mult_14_346 ;
wire Xd_0__inst_mult_14_348 ;
wire Xd_0__inst_mult_14_349 ;
wire Xd_0__inst_mult_14_350 ;
wire Xd_0__inst_mult_15_344 ;
wire Xd_0__inst_mult_15_345 ;
wire Xd_0__inst_mult_15_346 ;
wire Xd_0__inst_mult_15_348 ;
wire Xd_0__inst_mult_15_349 ;
wire Xd_0__inst_mult_15_350 ;
wire Xd_0__inst_mult_10_316 ;
wire Xd_0__inst_mult_10_317 ;
wire Xd_0__inst_mult_10_318 ;
wire Xd_0__inst_mult_10_320 ;
wire Xd_0__inst_mult_10_321 ;
wire Xd_0__inst_mult_10_322 ;
wire Xd_0__inst_mult_11_320 ;
wire Xd_0__inst_mult_11_321 ;
wire Xd_0__inst_mult_11_322 ;
wire Xd_0__inst_mult_11_324 ;
wire Xd_0__inst_mult_11_325 ;
wire Xd_0__inst_mult_11_326 ;
wire Xd_0__inst_mult_8_320 ;
wire Xd_0__inst_mult_8_321 ;
wire Xd_0__inst_mult_8_322 ;
wire Xd_0__inst_mult_8_324 ;
wire Xd_0__inst_mult_8_325 ;
wire Xd_0__inst_mult_8_326 ;
wire Xd_0__inst_mult_9_316 ;
wire Xd_0__inst_mult_9_317 ;
wire Xd_0__inst_mult_9_318 ;
wire Xd_0__inst_mult_9_320 ;
wire Xd_0__inst_mult_9_321 ;
wire Xd_0__inst_mult_9_322 ;
wire Xd_0__inst_mult_6_316 ;
wire Xd_0__inst_mult_6_317 ;
wire Xd_0__inst_mult_6_318 ;
wire Xd_0__inst_mult_6_320 ;
wire Xd_0__inst_mult_6_321 ;
wire Xd_0__inst_mult_6_322 ;
wire Xd_0__inst_mult_7_292 ;
wire Xd_0__inst_mult_7_293 ;
wire Xd_0__inst_mult_7_294 ;
wire Xd_0__inst_mult_7_296 ;
wire Xd_0__inst_mult_7_297 ;
wire Xd_0__inst_mult_7_298 ;
wire Xd_0__inst_mult_4_328 ;
wire Xd_0__inst_mult_4_329 ;
wire Xd_0__inst_mult_4_330 ;
wire Xd_0__inst_mult_4_332 ;
wire Xd_0__inst_mult_4_333 ;
wire Xd_0__inst_mult_4_334 ;
wire Xd_0__inst_mult_5_292 ;
wire Xd_0__inst_mult_5_293 ;
wire Xd_0__inst_mult_5_294 ;
wire Xd_0__inst_mult_5_296 ;
wire Xd_0__inst_mult_5_297 ;
wire Xd_0__inst_mult_5_298 ;
wire Xd_0__inst_mult_2_296 ;
wire Xd_0__inst_mult_2_297 ;
wire Xd_0__inst_mult_2_298 ;
wire Xd_0__inst_mult_2_300 ;
wire Xd_0__inst_mult_2_301 ;
wire Xd_0__inst_mult_2_302 ;
wire Xd_0__inst_mult_3_292 ;
wire Xd_0__inst_mult_3_293 ;
wire Xd_0__inst_mult_3_294 ;
wire Xd_0__inst_mult_3_296 ;
wire Xd_0__inst_mult_3_297 ;
wire Xd_0__inst_mult_3_298 ;
wire Xd_0__inst_mult_0_296 ;
wire Xd_0__inst_mult_0_297 ;
wire Xd_0__inst_mult_0_298 ;
wire Xd_0__inst_mult_0_300 ;
wire Xd_0__inst_mult_0_301 ;
wire Xd_0__inst_mult_0_302 ;
wire Xd_0__inst_mult_1_296 ;
wire Xd_0__inst_mult_1_297 ;
wire Xd_0__inst_mult_1_298 ;
wire Xd_0__inst_mult_1_300 ;
wire Xd_0__inst_mult_1_301 ;
wire Xd_0__inst_mult_1_302 ;
wire Xd_0__inst_mult_12_348 ;
wire Xd_0__inst_mult_12_349 ;
wire Xd_0__inst_mult_12_350 ;
wire Xd_0__inst_mult_12_352 ;
wire Xd_0__inst_mult_12_353 ;
wire Xd_0__inst_mult_12_354 ;
wire Xd_0__inst_mult_13_328 ;
wire Xd_0__inst_mult_13_329 ;
wire Xd_0__inst_mult_13_330 ;
wire Xd_0__inst_mult_13_332 ;
wire Xd_0__inst_mult_13_333 ;
wire Xd_0__inst_mult_13_334 ;
wire Xd_0__inst_mult_14_352 ;
wire Xd_0__inst_mult_14_353 ;
wire Xd_0__inst_mult_14_354 ;
wire Xd_0__inst_mult_14_356 ;
wire Xd_0__inst_mult_14_357 ;
wire Xd_0__inst_mult_14_358 ;
wire Xd_0__inst_mult_15_352 ;
wire Xd_0__inst_mult_15_353 ;
wire Xd_0__inst_mult_15_354 ;
wire Xd_0__inst_mult_15_356 ;
wire Xd_0__inst_mult_15_357 ;
wire Xd_0__inst_mult_15_358 ;
wire Xd_0__inst_mult_10_324 ;
wire Xd_0__inst_mult_10_325 ;
wire Xd_0__inst_mult_10_326 ;
wire Xd_0__inst_mult_10_328 ;
wire Xd_0__inst_mult_10_329 ;
wire Xd_0__inst_mult_10_330 ;
wire Xd_0__inst_mult_11_328 ;
wire Xd_0__inst_mult_11_329 ;
wire Xd_0__inst_mult_11_330 ;
wire Xd_0__inst_mult_11_332 ;
wire Xd_0__inst_mult_11_333 ;
wire Xd_0__inst_mult_11_334 ;
wire Xd_0__inst_mult_8_328 ;
wire Xd_0__inst_mult_8_329 ;
wire Xd_0__inst_mult_8_330 ;
wire Xd_0__inst_mult_8_332 ;
wire Xd_0__inst_mult_8_333 ;
wire Xd_0__inst_mult_8_334 ;
wire Xd_0__inst_mult_9_324 ;
wire Xd_0__inst_mult_9_325 ;
wire Xd_0__inst_mult_9_326 ;
wire Xd_0__inst_mult_9_328 ;
wire Xd_0__inst_mult_9_329 ;
wire Xd_0__inst_mult_9_330 ;
wire Xd_0__inst_mult_6_324 ;
wire Xd_0__inst_mult_6_325 ;
wire Xd_0__inst_mult_6_326 ;
wire Xd_0__inst_mult_6_328 ;
wire Xd_0__inst_mult_6_329 ;
wire Xd_0__inst_mult_6_330 ;
wire Xd_0__inst_mult_7_300 ;
wire Xd_0__inst_mult_7_301 ;
wire Xd_0__inst_mult_7_302 ;
wire Xd_0__inst_mult_7_304 ;
wire Xd_0__inst_mult_7_305 ;
wire Xd_0__inst_mult_7_306 ;
wire Xd_0__inst_mult_4_336 ;
wire Xd_0__inst_mult_4_337 ;
wire Xd_0__inst_mult_4_338 ;
wire Xd_0__inst_mult_4_340 ;
wire Xd_0__inst_mult_4_341 ;
wire Xd_0__inst_mult_4_342 ;
wire Xd_0__inst_mult_5_300 ;
wire Xd_0__inst_mult_5_301 ;
wire Xd_0__inst_mult_5_302 ;
wire Xd_0__inst_mult_5_304 ;
wire Xd_0__inst_mult_5_305 ;
wire Xd_0__inst_mult_5_306 ;
wire Xd_0__inst_mult_2_304 ;
wire Xd_0__inst_mult_2_305 ;
wire Xd_0__inst_mult_2_306 ;
wire Xd_0__inst_mult_2_308 ;
wire Xd_0__inst_mult_2_309 ;
wire Xd_0__inst_mult_2_310 ;
wire Xd_0__inst_mult_3_300 ;
wire Xd_0__inst_mult_3_301 ;
wire Xd_0__inst_mult_3_302 ;
wire Xd_0__inst_mult_3_304 ;
wire Xd_0__inst_mult_3_305 ;
wire Xd_0__inst_mult_3_306 ;
wire Xd_0__inst_mult_0_304 ;
wire Xd_0__inst_mult_0_305 ;
wire Xd_0__inst_mult_0_306 ;
wire Xd_0__inst_mult_0_308 ;
wire Xd_0__inst_mult_0_309 ;
wire Xd_0__inst_mult_0_310 ;
wire Xd_0__inst_mult_1_304 ;
wire Xd_0__inst_mult_1_305 ;
wire Xd_0__inst_mult_1_306 ;
wire Xd_0__inst_mult_1_308 ;
wire Xd_0__inst_mult_1_309 ;
wire Xd_0__inst_mult_1_310 ;
wire Xd_0__inst_mult_12_356 ;
wire Xd_0__inst_mult_12_357 ;
wire Xd_0__inst_mult_12_358 ;
wire Xd_0__inst_mult_12_360 ;
wire Xd_0__inst_mult_12_361 ;
wire Xd_0__inst_mult_12_362 ;
wire Xd_0__inst_mult_13_336 ;
wire Xd_0__inst_mult_13_337 ;
wire Xd_0__inst_mult_13_338 ;
wire Xd_0__inst_mult_13_340 ;
wire Xd_0__inst_mult_13_341 ;
wire Xd_0__inst_mult_13_342 ;
wire Xd_0__inst_mult_14_360 ;
wire Xd_0__inst_mult_14_361 ;
wire Xd_0__inst_mult_14_362 ;
wire Xd_0__inst_mult_15_360 ;
wire Xd_0__inst_mult_15_361 ;
wire Xd_0__inst_mult_15_362 ;
wire Xd_0__inst_mult_15_364 ;
wire Xd_0__inst_mult_15_365 ;
wire Xd_0__inst_mult_15_366 ;
wire Xd_0__inst_mult_10_332 ;
wire Xd_0__inst_mult_10_333 ;
wire Xd_0__inst_mult_10_334 ;
wire Xd_0__inst_mult_10_336 ;
wire Xd_0__inst_mult_10_337 ;
wire Xd_0__inst_mult_10_338 ;
wire Xd_0__inst_mult_11_336 ;
wire Xd_0__inst_mult_11_337 ;
wire Xd_0__inst_mult_11_338 ;
wire Xd_0__inst_mult_11_340 ;
wire Xd_0__inst_mult_11_341 ;
wire Xd_0__inst_mult_11_342 ;
wire Xd_0__inst_mult_8_336 ;
wire Xd_0__inst_mult_8_337 ;
wire Xd_0__inst_mult_8_338 ;
wire Xd_0__inst_mult_8_340 ;
wire Xd_0__inst_mult_8_341 ;
wire Xd_0__inst_mult_8_342 ;
wire Xd_0__inst_mult_9_332 ;
wire Xd_0__inst_mult_9_333 ;
wire Xd_0__inst_mult_9_334 ;
wire Xd_0__inst_mult_9_336 ;
wire Xd_0__inst_mult_9_337 ;
wire Xd_0__inst_mult_9_338 ;
wire Xd_0__inst_mult_6_332 ;
wire Xd_0__inst_mult_6_333 ;
wire Xd_0__inst_mult_6_334 ;
wire Xd_0__inst_mult_6_336 ;
wire Xd_0__inst_mult_6_337 ;
wire Xd_0__inst_mult_6_338 ;
wire Xd_0__inst_mult_7_308 ;
wire Xd_0__inst_mult_7_309 ;
wire Xd_0__inst_mult_7_310 ;
wire Xd_0__inst_mult_7_312 ;
wire Xd_0__inst_mult_7_313 ;
wire Xd_0__inst_mult_7_314 ;
wire Xd_0__inst_mult_4_344 ;
wire Xd_0__inst_mult_4_345 ;
wire Xd_0__inst_mult_4_346 ;
wire Xd_0__inst_mult_4_348 ;
wire Xd_0__inst_mult_4_349 ;
wire Xd_0__inst_mult_4_350 ;
wire Xd_0__inst_mult_5_308 ;
wire Xd_0__inst_mult_5_309 ;
wire Xd_0__inst_mult_5_310 ;
wire Xd_0__inst_mult_5_312 ;
wire Xd_0__inst_mult_5_313 ;
wire Xd_0__inst_mult_5_314 ;
wire Xd_0__inst_mult_2_312 ;
wire Xd_0__inst_mult_2_313 ;
wire Xd_0__inst_mult_2_314 ;
wire Xd_0__inst_mult_2_316 ;
wire Xd_0__inst_mult_2_317 ;
wire Xd_0__inst_mult_2_318 ;
wire Xd_0__inst_mult_3_308 ;
wire Xd_0__inst_mult_3_309 ;
wire Xd_0__inst_mult_3_310 ;
wire Xd_0__inst_mult_3_312 ;
wire Xd_0__inst_mult_3_313 ;
wire Xd_0__inst_mult_3_314 ;
wire Xd_0__inst_mult_0_312 ;
wire Xd_0__inst_mult_0_313 ;
wire Xd_0__inst_mult_0_314 ;
wire Xd_0__inst_mult_0_316 ;
wire Xd_0__inst_mult_0_317 ;
wire Xd_0__inst_mult_0_318 ;
wire Xd_0__inst_mult_1_312 ;
wire Xd_0__inst_mult_1_313 ;
wire Xd_0__inst_mult_1_314 ;
wire Xd_0__inst_mult_1_316 ;
wire Xd_0__inst_mult_1_317 ;
wire Xd_0__inst_mult_1_318 ;
wire Xd_0__inst_mult_12_364 ;
wire Xd_0__inst_mult_12_365 ;
wire Xd_0__inst_mult_12_366 ;
wire Xd_0__inst_mult_12_368 ;
wire Xd_0__inst_mult_12_369 ;
wire Xd_0__inst_mult_12_370 ;
wire Xd_0__inst_mult_13_344 ;
wire Xd_0__inst_mult_13_345 ;
wire Xd_0__inst_mult_13_346 ;
wire Xd_0__inst_mult_13_348 ;
wire Xd_0__inst_mult_13_349 ;
wire Xd_0__inst_mult_13_350 ;
wire Xd_0__inst_mult_14_364 ;
wire Xd_0__inst_mult_14_365 ;
wire Xd_0__inst_mult_14_366 ;
wire Xd_0__inst_mult_15_368 ;
wire Xd_0__inst_mult_15_369 ;
wire Xd_0__inst_mult_15_370 ;
wire Xd_0__inst_mult_15_372 ;
wire Xd_0__inst_mult_15_373 ;
wire Xd_0__inst_mult_15_374 ;
wire Xd_0__inst_mult_10_340 ;
wire Xd_0__inst_mult_10_341 ;
wire Xd_0__inst_mult_10_342 ;
wire Xd_0__inst_mult_10_344 ;
wire Xd_0__inst_mult_10_345 ;
wire Xd_0__inst_mult_10_346 ;
wire Xd_0__inst_mult_11_344 ;
wire Xd_0__inst_mult_11_345 ;
wire Xd_0__inst_mult_11_346 ;
wire Xd_0__inst_mult_11_348 ;
wire Xd_0__inst_mult_11_349 ;
wire Xd_0__inst_mult_11_350 ;
wire Xd_0__inst_mult_8_344 ;
wire Xd_0__inst_mult_8_345 ;
wire Xd_0__inst_mult_8_346 ;
wire Xd_0__inst_mult_8_348 ;
wire Xd_0__inst_mult_8_349 ;
wire Xd_0__inst_mult_8_350 ;
wire Xd_0__inst_mult_9_340 ;
wire Xd_0__inst_mult_9_341 ;
wire Xd_0__inst_mult_9_342 ;
wire Xd_0__inst_mult_9_344 ;
wire Xd_0__inst_mult_9_345 ;
wire Xd_0__inst_mult_9_346 ;
wire Xd_0__inst_mult_6_340 ;
wire Xd_0__inst_mult_6_341 ;
wire Xd_0__inst_mult_6_342 ;
wire Xd_0__inst_mult_6_344 ;
wire Xd_0__inst_mult_6_345 ;
wire Xd_0__inst_mult_6_346 ;
wire Xd_0__inst_mult_7_316 ;
wire Xd_0__inst_mult_7_317 ;
wire Xd_0__inst_mult_7_318 ;
wire Xd_0__inst_mult_7_320 ;
wire Xd_0__inst_mult_7_321 ;
wire Xd_0__inst_mult_7_322 ;
wire Xd_0__inst_mult_4_352 ;
wire Xd_0__inst_mult_4_353 ;
wire Xd_0__inst_mult_4_354 ;
wire Xd_0__inst_mult_4_356 ;
wire Xd_0__inst_mult_4_357 ;
wire Xd_0__inst_mult_4_358 ;
wire Xd_0__inst_mult_5_316 ;
wire Xd_0__inst_mult_5_317 ;
wire Xd_0__inst_mult_5_318 ;
wire Xd_0__inst_mult_5_320 ;
wire Xd_0__inst_mult_5_321 ;
wire Xd_0__inst_mult_5_322 ;
wire Xd_0__inst_mult_2_320 ;
wire Xd_0__inst_mult_2_321 ;
wire Xd_0__inst_mult_2_322 ;
wire Xd_0__inst_mult_2_324 ;
wire Xd_0__inst_mult_2_325 ;
wire Xd_0__inst_mult_2_326 ;
wire Xd_0__inst_mult_3_316 ;
wire Xd_0__inst_mult_3_317 ;
wire Xd_0__inst_mult_3_318 ;
wire Xd_0__inst_mult_3_320 ;
wire Xd_0__inst_mult_3_321 ;
wire Xd_0__inst_mult_3_322 ;
wire Xd_0__inst_mult_0_320 ;
wire Xd_0__inst_mult_0_321 ;
wire Xd_0__inst_mult_0_322 ;
wire Xd_0__inst_mult_0_324 ;
wire Xd_0__inst_mult_0_325 ;
wire Xd_0__inst_mult_0_326 ;
wire Xd_0__inst_mult_1_320 ;
wire Xd_0__inst_mult_1_321 ;
wire Xd_0__inst_mult_1_322 ;
wire Xd_0__inst_mult_1_324 ;
wire Xd_0__inst_mult_1_325 ;
wire Xd_0__inst_mult_1_326 ;
wire Xd_0__inst_mult_12_372 ;
wire Xd_0__inst_mult_12_373 ;
wire Xd_0__inst_mult_12_374 ;
wire Xd_0__inst_mult_13_352 ;
wire Xd_0__inst_mult_13_353 ;
wire Xd_0__inst_mult_13_354 ;
wire Xd_0__inst_mult_14_368 ;
wire Xd_0__inst_mult_14_369 ;
wire Xd_0__inst_mult_14_370 ;
wire Xd_0__inst_mult_15_376 ;
wire Xd_0__inst_mult_15_377 ;
wire Xd_0__inst_mult_15_378 ;
wire Xd_0__inst_mult_10_348 ;
wire Xd_0__inst_mult_10_349 ;
wire Xd_0__inst_mult_10_350 ;
wire Xd_0__inst_mult_11_352 ;
wire Xd_0__inst_mult_11_353 ;
wire Xd_0__inst_mult_11_354 ;
wire Xd_0__inst_mult_8_352 ;
wire Xd_0__inst_mult_8_353 ;
wire Xd_0__inst_mult_8_354 ;
wire Xd_0__inst_mult_9_348 ;
wire Xd_0__inst_mult_9_349 ;
wire Xd_0__inst_mult_9_350 ;
wire Xd_0__inst_mult_6_348 ;
wire Xd_0__inst_mult_6_349 ;
wire Xd_0__inst_mult_6_350 ;
wire Xd_0__inst_mult_7_324 ;
wire Xd_0__inst_mult_7_325 ;
wire Xd_0__inst_mult_7_326 ;
wire Xd_0__inst_mult_7_328 ;
wire Xd_0__inst_mult_7_329 ;
wire Xd_0__inst_mult_7_330 ;
wire Xd_0__inst_mult_4_360 ;
wire Xd_0__inst_mult_4_361 ;
wire Xd_0__inst_mult_4_362 ;
wire Xd_0__inst_mult_4_364 ;
wire Xd_0__inst_mult_4_365 ;
wire Xd_0__inst_mult_4_366 ;
wire Xd_0__inst_mult_5_324 ;
wire Xd_0__inst_mult_5_325 ;
wire Xd_0__inst_mult_5_326 ;
wire Xd_0__inst_mult_5_328 ;
wire Xd_0__inst_mult_5_329 ;
wire Xd_0__inst_mult_5_330 ;
wire Xd_0__inst_mult_2_328 ;
wire Xd_0__inst_mult_2_329 ;
wire Xd_0__inst_mult_2_330 ;
wire Xd_0__inst_mult_2_332 ;
wire Xd_0__inst_mult_2_333 ;
wire Xd_0__inst_mult_2_334 ;
wire Xd_0__inst_mult_3_324 ;
wire Xd_0__inst_mult_3_325 ;
wire Xd_0__inst_mult_3_326 ;
wire Xd_0__inst_mult_3_328 ;
wire Xd_0__inst_mult_3_329 ;
wire Xd_0__inst_mult_3_330 ;
wire Xd_0__inst_mult_0_328 ;
wire Xd_0__inst_mult_0_329 ;
wire Xd_0__inst_mult_0_330 ;
wire Xd_0__inst_mult_0_332 ;
wire Xd_0__inst_mult_0_333 ;
wire Xd_0__inst_mult_0_334 ;
wire Xd_0__inst_mult_1_328 ;
wire Xd_0__inst_mult_1_329 ;
wire Xd_0__inst_mult_1_330 ;
wire Xd_0__inst_mult_1_332 ;
wire Xd_0__inst_mult_1_333 ;
wire Xd_0__inst_mult_1_334 ;
wire Xd_0__inst_mult_12_376 ;
wire Xd_0__inst_mult_12_377 ;
wire Xd_0__inst_mult_12_378 ;
wire Xd_0__inst_mult_13_356 ;
wire Xd_0__inst_mult_13_357 ;
wire Xd_0__inst_mult_13_358 ;
wire Xd_0__inst_mult_14_372 ;
wire Xd_0__inst_mult_14_373 ;
wire Xd_0__inst_mult_14_374 ;
wire Xd_0__inst_mult_15_380 ;
wire Xd_0__inst_mult_15_381 ;
wire Xd_0__inst_mult_15_382 ;
wire Xd_0__inst_mult_10_352 ;
wire Xd_0__inst_mult_10_353 ;
wire Xd_0__inst_mult_10_354 ;
wire Xd_0__inst_mult_11_356 ;
wire Xd_0__inst_mult_11_357 ;
wire Xd_0__inst_mult_11_358 ;
wire Xd_0__inst_mult_8_356 ;
wire Xd_0__inst_mult_8_357 ;
wire Xd_0__inst_mult_8_358 ;
wire Xd_0__inst_mult_9_352 ;
wire Xd_0__inst_mult_9_353 ;
wire Xd_0__inst_mult_9_354 ;
wire Xd_0__inst_mult_6_352 ;
wire Xd_0__inst_mult_6_353 ;
wire Xd_0__inst_mult_6_354 ;
wire Xd_0__inst_mult_7_332 ;
wire Xd_0__inst_mult_7_333 ;
wire Xd_0__inst_mult_7_334 ;
wire Xd_0__inst_mult_7_336 ;
wire Xd_0__inst_mult_7_337 ;
wire Xd_0__inst_mult_7_338 ;
wire Xd_0__inst_mult_4_368 ;
wire Xd_0__inst_mult_4_369 ;
wire Xd_0__inst_mult_4_370 ;
wire Xd_0__inst_mult_4_372 ;
wire Xd_0__inst_mult_4_373 ;
wire Xd_0__inst_mult_4_374 ;
wire Xd_0__inst_mult_5_332 ;
wire Xd_0__inst_mult_5_333 ;
wire Xd_0__inst_mult_5_334 ;
wire Xd_0__inst_mult_5_336 ;
wire Xd_0__inst_mult_5_337 ;
wire Xd_0__inst_mult_5_338 ;
wire Xd_0__inst_mult_2_336 ;
wire Xd_0__inst_mult_2_337 ;
wire Xd_0__inst_mult_2_338 ;
wire Xd_0__inst_mult_2_340 ;
wire Xd_0__inst_mult_2_341 ;
wire Xd_0__inst_mult_2_342 ;
wire Xd_0__inst_mult_3_332 ;
wire Xd_0__inst_mult_3_333 ;
wire Xd_0__inst_mult_3_334 ;
wire Xd_0__inst_mult_3_336 ;
wire Xd_0__inst_mult_3_337 ;
wire Xd_0__inst_mult_3_338 ;
wire Xd_0__inst_mult_0_336 ;
wire Xd_0__inst_mult_0_337 ;
wire Xd_0__inst_mult_0_338 ;
wire Xd_0__inst_mult_0_340 ;
wire Xd_0__inst_mult_0_341 ;
wire Xd_0__inst_mult_0_342 ;
wire Xd_0__inst_mult_1_336 ;
wire Xd_0__inst_mult_1_337 ;
wire Xd_0__inst_mult_1_338 ;
wire Xd_0__inst_mult_1_340 ;
wire Xd_0__inst_mult_1_341 ;
wire Xd_0__inst_mult_1_342 ;
wire Xd_0__inst_mult_12_380 ;
wire Xd_0__inst_mult_12_381 ;
wire Xd_0__inst_mult_12_382 ;
wire Xd_0__inst_mult_13_360 ;
wire Xd_0__inst_mult_13_361 ;
wire Xd_0__inst_mult_13_362 ;
wire Xd_0__inst_mult_14_376 ;
wire Xd_0__inst_mult_14_377 ;
wire Xd_0__inst_mult_14_378 ;
wire Xd_0__inst_mult_15_384 ;
wire Xd_0__inst_mult_15_385 ;
wire Xd_0__inst_mult_15_386 ;
wire Xd_0__inst_mult_10_356 ;
wire Xd_0__inst_mult_10_357 ;
wire Xd_0__inst_mult_10_358 ;
wire Xd_0__inst_mult_11_360 ;
wire Xd_0__inst_mult_11_361 ;
wire Xd_0__inst_mult_11_362 ;
wire Xd_0__inst_mult_8_360 ;
wire Xd_0__inst_mult_8_361 ;
wire Xd_0__inst_mult_8_362 ;
wire Xd_0__inst_mult_9_356 ;
wire Xd_0__inst_mult_9_357 ;
wire Xd_0__inst_mult_9_358 ;
wire Xd_0__inst_mult_6_356 ;
wire Xd_0__inst_mult_6_357 ;
wire Xd_0__inst_mult_6_358 ;
wire Xd_0__inst_mult_7_340 ;
wire Xd_0__inst_mult_7_341 ;
wire Xd_0__inst_mult_7_342 ;
wire Xd_0__inst_mult_7_344 ;
wire Xd_0__inst_mult_7_345 ;
wire Xd_0__inst_mult_7_346 ;
wire Xd_0__inst_mult_4_376 ;
wire Xd_0__inst_mult_4_377 ;
wire Xd_0__inst_mult_4_378 ;
wire Xd_0__inst_mult_4_380 ;
wire Xd_0__inst_mult_4_381 ;
wire Xd_0__inst_mult_4_382 ;
wire Xd_0__inst_mult_5_340 ;
wire Xd_0__inst_mult_5_341 ;
wire Xd_0__inst_mult_5_342 ;
wire Xd_0__inst_mult_5_344 ;
wire Xd_0__inst_mult_5_345 ;
wire Xd_0__inst_mult_5_346 ;
wire Xd_0__inst_mult_2_344 ;
wire Xd_0__inst_mult_2_345 ;
wire Xd_0__inst_mult_2_346 ;
wire Xd_0__inst_mult_2_348 ;
wire Xd_0__inst_mult_2_349 ;
wire Xd_0__inst_mult_2_350 ;
wire Xd_0__inst_mult_3_340 ;
wire Xd_0__inst_mult_3_341 ;
wire Xd_0__inst_mult_3_342 ;
wire Xd_0__inst_mult_3_344 ;
wire Xd_0__inst_mult_3_345 ;
wire Xd_0__inst_mult_3_346 ;
wire Xd_0__inst_mult_0_344 ;
wire Xd_0__inst_mult_0_345 ;
wire Xd_0__inst_mult_0_346 ;
wire Xd_0__inst_mult_0_348 ;
wire Xd_0__inst_mult_0_349 ;
wire Xd_0__inst_mult_0_350 ;
wire Xd_0__inst_mult_1_344 ;
wire Xd_0__inst_mult_1_345 ;
wire Xd_0__inst_mult_1_346 ;
wire Xd_0__inst_mult_1_348 ;
wire Xd_0__inst_mult_1_349 ;
wire Xd_0__inst_mult_1_350 ;
wire Xd_0__inst_mult_12_384 ;
wire Xd_0__inst_mult_12_385 ;
wire Xd_0__inst_mult_12_386 ;
wire Xd_0__inst_mult_13_364 ;
wire Xd_0__inst_mult_13_365 ;
wire Xd_0__inst_mult_13_366 ;
wire Xd_0__inst_mult_14_380 ;
wire Xd_0__inst_mult_14_381 ;
wire Xd_0__inst_mult_14_382 ;
wire Xd_0__inst_mult_15_388 ;
wire Xd_0__inst_mult_15_389 ;
wire Xd_0__inst_mult_15_390 ;
wire Xd_0__inst_mult_10_360 ;
wire Xd_0__inst_mult_10_361 ;
wire Xd_0__inst_mult_10_362 ;
wire Xd_0__inst_mult_11_364 ;
wire Xd_0__inst_mult_11_365 ;
wire Xd_0__inst_mult_11_366 ;
wire Xd_0__inst_mult_8_364 ;
wire Xd_0__inst_mult_8_365 ;
wire Xd_0__inst_mult_8_366 ;
wire Xd_0__inst_mult_9_360 ;
wire Xd_0__inst_mult_9_361 ;
wire Xd_0__inst_mult_9_362 ;
wire Xd_0__inst_mult_6_360 ;
wire Xd_0__inst_mult_6_361 ;
wire Xd_0__inst_mult_6_362 ;
wire Xd_0__inst_mult_7_348 ;
wire Xd_0__inst_mult_7_352 ;
wire Xd_0__inst_mult_7_353 ;
wire Xd_0__inst_mult_7_354 ;
wire Xd_0__inst_mult_4_384 ;
wire Xd_0__inst_mult_4_388 ;
wire Xd_0__inst_mult_4_389 ;
wire Xd_0__inst_mult_4_390 ;
wire Xd_0__inst_mult_5_348 ;
wire Xd_0__inst_mult_5_352 ;
wire Xd_0__inst_mult_5_353 ;
wire Xd_0__inst_mult_5_354 ;
wire Xd_0__inst_mult_2_352 ;
wire Xd_0__inst_mult_2_356 ;
wire Xd_0__inst_mult_2_357 ;
wire Xd_0__inst_mult_2_358 ;
wire Xd_0__inst_mult_3_348 ;
wire Xd_0__inst_mult_3_352 ;
wire Xd_0__inst_mult_3_353 ;
wire Xd_0__inst_mult_3_354 ;
wire Xd_0__inst_mult_0_352 ;
wire Xd_0__inst_mult_0_356 ;
wire Xd_0__inst_mult_0_357 ;
wire Xd_0__inst_mult_0_358 ;
wire Xd_0__inst_mult_1_352 ;
wire Xd_0__inst_mult_1_356 ;
wire Xd_0__inst_mult_1_357 ;
wire Xd_0__inst_mult_1_358 ;
wire Xd_0__inst_mult_12_388 ;
wire Xd_0__inst_mult_12_389 ;
wire Xd_0__inst_mult_12_390 ;
wire Xd_0__inst_mult_12_47_sumout ;
wire Xd_0__inst_mult_12_48 ;
wire Xd_0__inst_mult_12_49 ;
wire Xd_0__inst_mult_13_368 ;
wire Xd_0__inst_mult_13_369 ;
wire Xd_0__inst_mult_13_370 ;
wire Xd_0__inst_mult_13_43_sumout ;
wire Xd_0__inst_mult_13_44 ;
wire Xd_0__inst_mult_13_45 ;
wire Xd_0__inst_mult_14_384 ;
wire Xd_0__inst_mult_14_385 ;
wire Xd_0__inst_mult_14_386 ;
wire Xd_0__inst_mult_15_392 ;
wire Xd_0__inst_mult_15_393 ;
wire Xd_0__inst_mult_15_394 ;
wire Xd_0__inst_mult_15_47_sumout ;
wire Xd_0__inst_mult_15_48 ;
wire Xd_0__inst_mult_15_49 ;
wire Xd_0__inst_mult_10_364 ;
wire Xd_0__inst_mult_10_365 ;
wire Xd_0__inst_mult_10_366 ;
wire Xd_0__inst_mult_0_360 ;
wire Xd_0__inst_mult_0_361 ;
wire Xd_0__inst_mult_0_362 ;
wire Xd_0__inst_mult_11_368 ;
wire Xd_0__inst_mult_11_369 ;
wire Xd_0__inst_mult_11_370 ;
wire Xd_0__inst_mult_11_39_sumout ;
wire Xd_0__inst_mult_11_40 ;
wire Xd_0__inst_mult_11_41 ;
wire Xd_0__inst_mult_8_368 ;
wire Xd_0__inst_mult_8_369 ;
wire Xd_0__inst_mult_8_370 ;
wire Xd_0__inst_mult_8_47_sumout ;
wire Xd_0__inst_mult_8_48 ;
wire Xd_0__inst_mult_8_49 ;
wire Xd_0__inst_mult_9_364 ;
wire Xd_0__inst_mult_9_365 ;
wire Xd_0__inst_mult_9_366 ;
wire Xd_0__inst_mult_9_39_sumout ;
wire Xd_0__inst_mult_9_40 ;
wire Xd_0__inst_mult_9_41 ;
wire Xd_0__inst_mult_6_364 ;
wire Xd_0__inst_mult_6_365 ;
wire Xd_0__inst_mult_6_366 ;
wire Xd_0__inst_mult_6_43_sumout ;
wire Xd_0__inst_mult_6_44 ;
wire Xd_0__inst_mult_6_45 ;
wire Xd_0__inst_mult_7_356 ;
wire Xd_0__inst_mult_7_357 ;
wire Xd_0__inst_mult_7_358 ;
wire Xd_0__inst_mult_1_360 ;
wire Xd_0__inst_mult_1_361 ;
wire Xd_0__inst_mult_1_362 ;
wire Xd_0__inst_mult_4_392 ;
wire Xd_0__inst_mult_4_393 ;
wire Xd_0__inst_mult_4_394 ;
wire Xd_0__inst_mult_4_39_sumout ;
wire Xd_0__inst_mult_4_40 ;
wire Xd_0__inst_mult_4_41 ;
wire Xd_0__inst_mult_5_356 ;
wire Xd_0__inst_mult_5_357 ;
wire Xd_0__inst_mult_5_358 ;
wire Xd_0__inst_mult_5_43_sumout ;
wire Xd_0__inst_mult_5_44 ;
wire Xd_0__inst_mult_5_45 ;
wire Xd_0__inst_mult_2_360 ;
wire Xd_0__inst_mult_2_361 ;
wire Xd_0__inst_mult_2_362 ;
wire Xd_0__inst_mult_2_43_sumout ;
wire Xd_0__inst_mult_2_44 ;
wire Xd_0__inst_mult_2_45 ;
wire Xd_0__inst_mult_3_356 ;
wire Xd_0__inst_mult_3_357 ;
wire Xd_0__inst_mult_3_358 ;
wire Xd_0__inst_mult_3_47_sumout ;
wire Xd_0__inst_mult_3_48 ;
wire Xd_0__inst_mult_3_49 ;
wire Xd_0__inst_mult_0_364 ;
wire Xd_0__inst_mult_0_365 ;
wire Xd_0__inst_mult_0_366 ;
wire Xd_0__inst_mult_0_39_sumout ;
wire Xd_0__inst_mult_0_40 ;
wire Xd_0__inst_mult_0_41 ;
wire Xd_0__inst_mult_1_364 ;
wire Xd_0__inst_mult_1_365 ;
wire Xd_0__inst_mult_1_366 ;
wire Xd_0__inst_mult_1_43_sumout ;
wire Xd_0__inst_mult_1_44 ;
wire Xd_0__inst_mult_1_45 ;
wire Xd_0__inst_mult_12_392 ;
wire Xd_0__inst_mult_12_393 ;
wire Xd_0__inst_mult_12_394 ;
wire Xd_0__inst_mult_12_51_sumout ;
wire Xd_0__inst_mult_12_52 ;
wire Xd_0__inst_mult_12_53 ;
wire Xd_0__inst_mult_13_372 ;
wire Xd_0__inst_mult_13_373 ;
wire Xd_0__inst_mult_13_374 ;
wire Xd_0__inst_mult_13_47_sumout ;
wire Xd_0__inst_mult_13_48 ;
wire Xd_0__inst_mult_13_49 ;
wire Xd_0__inst_mult_14_388 ;
wire Xd_0__inst_mult_14_389 ;
wire Xd_0__inst_mult_14_390 ;
wire Xd_0__inst_mult_14_55_sumout ;
wire Xd_0__inst_mult_14_56 ;
wire Xd_0__inst_mult_14_57 ;
wire Xd_0__inst_mult_15_396 ;
wire Xd_0__inst_mult_15_397 ;
wire Xd_0__inst_mult_15_398 ;
wire Xd_0__inst_mult_15_51_sumout ;
wire Xd_0__inst_mult_15_52 ;
wire Xd_0__inst_mult_15_53 ;
wire Xd_0__inst_mult_10_368 ;
wire Xd_0__inst_mult_10_369 ;
wire Xd_0__inst_mult_10_370 ;
wire Xd_0__inst_mult_10_43_sumout ;
wire Xd_0__inst_mult_10_44 ;
wire Xd_0__inst_mult_10_45 ;
wire Xd_0__inst_mult_11_372 ;
wire Xd_0__inst_mult_11_373 ;
wire Xd_0__inst_mult_11_374 ;
wire Xd_0__inst_mult_11_43_sumout ;
wire Xd_0__inst_mult_11_44 ;
wire Xd_0__inst_mult_11_45 ;
wire Xd_0__inst_mult_8_372 ;
wire Xd_0__inst_mult_8_373 ;
wire Xd_0__inst_mult_8_374 ;
wire Xd_0__inst_mult_8_51_sumout ;
wire Xd_0__inst_mult_8_52 ;
wire Xd_0__inst_mult_8_53 ;
wire Xd_0__inst_mult_9_368 ;
wire Xd_0__inst_mult_9_369 ;
wire Xd_0__inst_mult_9_370 ;
wire Xd_0__inst_mult_6_368 ;
wire Xd_0__inst_mult_6_369 ;
wire Xd_0__inst_mult_6_370 ;
wire Xd_0__inst_mult_6_47_sumout ;
wire Xd_0__inst_mult_6_48 ;
wire Xd_0__inst_mult_6_49 ;
wire Xd_0__inst_mult_7_360 ;
wire Xd_0__inst_mult_7_361 ;
wire Xd_0__inst_mult_7_362 ;
wire Xd_0__inst_mult_7_39_sumout ;
wire Xd_0__inst_mult_7_40 ;
wire Xd_0__inst_mult_7_41 ;
wire Xd_0__inst_mult_4_396 ;
wire Xd_0__inst_mult_4_397 ;
wire Xd_0__inst_mult_4_398 ;
wire Xd_0__inst_mult_4_43_sumout ;
wire Xd_0__inst_mult_4_44 ;
wire Xd_0__inst_mult_4_45 ;
wire Xd_0__inst_mult_5_360 ;
wire Xd_0__inst_mult_5_361 ;
wire Xd_0__inst_mult_5_362 ;
wire Xd_0__inst_mult_5_47_sumout ;
wire Xd_0__inst_mult_5_48 ;
wire Xd_0__inst_mult_5_49 ;
wire Xd_0__inst_mult_2_364 ;
wire Xd_0__inst_mult_2_365 ;
wire Xd_0__inst_mult_2_366 ;
wire Xd_0__inst_mult_2_47_sumout ;
wire Xd_0__inst_mult_2_48 ;
wire Xd_0__inst_mult_2_49 ;
wire Xd_0__inst_mult_3_360 ;
wire Xd_0__inst_mult_3_361 ;
wire Xd_0__inst_mult_3_362 ;
wire Xd_0__inst_mult_3_51_sumout ;
wire Xd_0__inst_mult_3_52 ;
wire Xd_0__inst_mult_3_53 ;
wire Xd_0__inst_mult_0_368 ;
wire Xd_0__inst_mult_0_369 ;
wire Xd_0__inst_mult_0_370 ;
wire Xd_0__inst_mult_0_43_sumout ;
wire Xd_0__inst_mult_0_44 ;
wire Xd_0__inst_mult_0_45 ;
wire Xd_0__inst_mult_1_368 ;
wire Xd_0__inst_mult_1_369 ;
wire Xd_0__inst_mult_1_370 ;
wire Xd_0__inst_mult_1_47_sumout ;
wire Xd_0__inst_mult_1_48 ;
wire Xd_0__inst_mult_1_49 ;
wire Xd_0__inst_mult_12_396 ;
wire Xd_0__inst_mult_12_397 ;
wire Xd_0__inst_mult_12_398 ;
wire Xd_0__inst_mult_12_55_sumout ;
wire Xd_0__inst_mult_12_56 ;
wire Xd_0__inst_mult_12_57 ;
wire Xd_0__inst_mult_13_376 ;
wire Xd_0__inst_mult_13_377 ;
wire Xd_0__inst_mult_13_378 ;
wire Xd_0__inst_mult_13_51_sumout ;
wire Xd_0__inst_mult_13_52 ;
wire Xd_0__inst_mult_13_53 ;
wire Xd_0__inst_mult_14_392 ;
wire Xd_0__inst_mult_14_393 ;
wire Xd_0__inst_mult_14_394 ;
wire Xd_0__inst_mult_14_59_sumout ;
wire Xd_0__inst_mult_14_60 ;
wire Xd_0__inst_mult_14_61 ;
wire Xd_0__inst_mult_15_400 ;
wire Xd_0__inst_mult_15_401 ;
wire Xd_0__inst_mult_15_402 ;
wire Xd_0__inst_mult_15_55_sumout ;
wire Xd_0__inst_mult_15_56 ;
wire Xd_0__inst_mult_15_57 ;
wire Xd_0__inst_mult_10_372 ;
wire Xd_0__inst_mult_10_373 ;
wire Xd_0__inst_mult_10_374 ;
wire Xd_0__inst_mult_10_47_sumout ;
wire Xd_0__inst_mult_10_48 ;
wire Xd_0__inst_mult_10_49 ;
wire Xd_0__inst_mult_11_376 ;
wire Xd_0__inst_mult_11_377 ;
wire Xd_0__inst_mult_11_378 ;
wire Xd_0__inst_mult_11_47_sumout ;
wire Xd_0__inst_mult_11_48 ;
wire Xd_0__inst_mult_11_49 ;
wire Xd_0__inst_mult_8_376 ;
wire Xd_0__inst_mult_8_377 ;
wire Xd_0__inst_mult_8_378 ;
wire Xd_0__inst_mult_8_55_sumout ;
wire Xd_0__inst_mult_8_56 ;
wire Xd_0__inst_mult_8_57 ;
wire Xd_0__inst_mult_9_372 ;
wire Xd_0__inst_mult_9_373 ;
wire Xd_0__inst_mult_9_374 ;
wire Xd_0__inst_mult_9_43_sumout ;
wire Xd_0__inst_mult_9_44 ;
wire Xd_0__inst_mult_9_45 ;
wire Xd_0__inst_mult_6_372 ;
wire Xd_0__inst_mult_6_373 ;
wire Xd_0__inst_mult_6_374 ;
wire Xd_0__inst_mult_6_51_sumout ;
wire Xd_0__inst_mult_6_52 ;
wire Xd_0__inst_mult_6_53 ;
wire Xd_0__inst_mult_7_364 ;
wire Xd_0__inst_mult_7_365 ;
wire Xd_0__inst_mult_7_366 ;
wire Xd_0__inst_mult_7_43_sumout ;
wire Xd_0__inst_mult_7_44 ;
wire Xd_0__inst_mult_7_45 ;
wire Xd_0__inst_mult_4_400 ;
wire Xd_0__inst_mult_4_401 ;
wire Xd_0__inst_mult_4_402 ;
wire Xd_0__inst_mult_4_47_sumout ;
wire Xd_0__inst_mult_4_48 ;
wire Xd_0__inst_mult_4_49 ;
wire Xd_0__inst_mult_5_364 ;
wire Xd_0__inst_mult_5_365 ;
wire Xd_0__inst_mult_5_366 ;
wire Xd_0__inst_mult_5_51_sumout ;
wire Xd_0__inst_mult_5_52 ;
wire Xd_0__inst_mult_5_53 ;
wire Xd_0__inst_mult_2_368 ;
wire Xd_0__inst_mult_2_369 ;
wire Xd_0__inst_mult_2_370 ;
wire Xd_0__inst_mult_2_51_sumout ;
wire Xd_0__inst_mult_2_52 ;
wire Xd_0__inst_mult_2_53 ;
wire Xd_0__inst_mult_3_364 ;
wire Xd_0__inst_mult_3_365 ;
wire Xd_0__inst_mult_3_366 ;
wire Xd_0__inst_mult_3_55_sumout ;
wire Xd_0__inst_mult_3_56 ;
wire Xd_0__inst_mult_3_57 ;
wire Xd_0__inst_mult_0_372 ;
wire Xd_0__inst_mult_0_373 ;
wire Xd_0__inst_mult_0_374 ;
wire Xd_0__inst_mult_0_47_sumout ;
wire Xd_0__inst_mult_0_48 ;
wire Xd_0__inst_mult_0_49 ;
wire Xd_0__inst_mult_1_372 ;
wire Xd_0__inst_mult_1_373 ;
wire Xd_0__inst_mult_1_374 ;
wire Xd_0__inst_mult_1_51_sumout ;
wire Xd_0__inst_mult_1_52 ;
wire Xd_0__inst_mult_1_53 ;
wire Xd_0__inst_mult_12_400 ;
wire Xd_0__inst_mult_12_401 ;
wire Xd_0__inst_mult_12_402 ;
wire Xd_0__inst_mult_12_59_sumout ;
wire Xd_0__inst_mult_12_60 ;
wire Xd_0__inst_mult_12_61 ;
wire Xd_0__inst_mult_13_380 ;
wire Xd_0__inst_mult_13_381 ;
wire Xd_0__inst_mult_13_382 ;
wire Xd_0__inst_mult_13_55_sumout ;
wire Xd_0__inst_mult_13_56 ;
wire Xd_0__inst_mult_13_57 ;
wire Xd_0__inst_mult_14_396 ;
wire Xd_0__inst_mult_14_397 ;
wire Xd_0__inst_mult_14_398 ;
wire Xd_0__inst_mult_14_63_sumout ;
wire Xd_0__inst_mult_14_64 ;
wire Xd_0__inst_mult_14_65 ;
wire Xd_0__inst_mult_15_404 ;
wire Xd_0__inst_mult_15_405 ;
wire Xd_0__inst_mult_15_406 ;
wire Xd_0__inst_mult_15_59_sumout ;
wire Xd_0__inst_mult_15_60 ;
wire Xd_0__inst_mult_15_61 ;
wire Xd_0__inst_mult_10_376 ;
wire Xd_0__inst_mult_10_377 ;
wire Xd_0__inst_mult_10_378 ;
wire Xd_0__inst_mult_10_51_sumout ;
wire Xd_0__inst_mult_10_52 ;
wire Xd_0__inst_mult_10_53 ;
wire Xd_0__inst_mult_11_380 ;
wire Xd_0__inst_mult_11_381 ;
wire Xd_0__inst_mult_11_382 ;
wire Xd_0__inst_mult_11_51_sumout ;
wire Xd_0__inst_mult_11_52 ;
wire Xd_0__inst_mult_11_53 ;
wire Xd_0__inst_mult_8_380 ;
wire Xd_0__inst_mult_8_381 ;
wire Xd_0__inst_mult_8_382 ;
wire Xd_0__inst_mult_8_59_sumout ;
wire Xd_0__inst_mult_8_60 ;
wire Xd_0__inst_mult_8_61 ;
wire Xd_0__inst_mult_9_376 ;
wire Xd_0__inst_mult_9_377 ;
wire Xd_0__inst_mult_9_378 ;
wire Xd_0__inst_mult_9_47_sumout ;
wire Xd_0__inst_mult_9_48 ;
wire Xd_0__inst_mult_9_49 ;
wire Xd_0__inst_mult_6_376 ;
wire Xd_0__inst_mult_6_377 ;
wire Xd_0__inst_mult_6_378 ;
wire Xd_0__inst_mult_6_55_sumout ;
wire Xd_0__inst_mult_6_56 ;
wire Xd_0__inst_mult_6_57 ;
wire Xd_0__inst_mult_7_368 ;
wire Xd_0__inst_mult_7_369 ;
wire Xd_0__inst_mult_7_370 ;
wire Xd_0__inst_mult_7_47_sumout ;
wire Xd_0__inst_mult_7_48 ;
wire Xd_0__inst_mult_7_49 ;
wire Xd_0__inst_mult_4_404 ;
wire Xd_0__inst_mult_4_405 ;
wire Xd_0__inst_mult_4_406 ;
wire Xd_0__inst_mult_4_51_sumout ;
wire Xd_0__inst_mult_4_52 ;
wire Xd_0__inst_mult_4_53 ;
wire Xd_0__inst_mult_5_368 ;
wire Xd_0__inst_mult_5_369 ;
wire Xd_0__inst_mult_5_370 ;
wire Xd_0__inst_mult_5_55_sumout ;
wire Xd_0__inst_mult_5_56 ;
wire Xd_0__inst_mult_5_57 ;
wire Xd_0__inst_mult_2_372 ;
wire Xd_0__inst_mult_2_373 ;
wire Xd_0__inst_mult_2_374 ;
wire Xd_0__inst_mult_2_55_sumout ;
wire Xd_0__inst_mult_2_56 ;
wire Xd_0__inst_mult_2_57 ;
wire Xd_0__inst_mult_3_368 ;
wire Xd_0__inst_mult_3_369 ;
wire Xd_0__inst_mult_3_370 ;
wire Xd_0__inst_mult_3_59_sumout ;
wire Xd_0__inst_mult_3_60 ;
wire Xd_0__inst_mult_3_61 ;
wire Xd_0__inst_mult_0_376 ;
wire Xd_0__inst_mult_0_377 ;
wire Xd_0__inst_mult_0_378 ;
wire Xd_0__inst_mult_0_51_sumout ;
wire Xd_0__inst_mult_0_52 ;
wire Xd_0__inst_mult_0_53 ;
wire Xd_0__inst_mult_1_376 ;
wire Xd_0__inst_mult_1_377 ;
wire Xd_0__inst_mult_1_378 ;
wire Xd_0__inst_mult_1_55_sumout ;
wire Xd_0__inst_mult_1_56 ;
wire Xd_0__inst_mult_1_57 ;
wire Xd_0__inst_mult_12_404 ;
wire Xd_0__inst_mult_13_384 ;
wire Xd_0__inst_mult_13_59_sumout ;
wire Xd_0__inst_mult_13_60 ;
wire Xd_0__inst_mult_13_61 ;
wire Xd_0__inst_mult_14_400 ;
wire Xd_0__inst_mult_15_408 ;
wire Xd_0__inst_mult_10_380 ;
wire Xd_0__inst_mult_10_55_sumout ;
wire Xd_0__inst_mult_10_56 ;
wire Xd_0__inst_mult_10_57 ;
wire Xd_0__inst_mult_11_384 ;
wire Xd_0__inst_mult_8_384 ;
wire Xd_0__inst_mult_9_380 ;
wire Xd_0__inst_mult_9_51_sumout ;
wire Xd_0__inst_mult_9_52 ;
wire Xd_0__inst_mult_9_53 ;
wire Xd_0__inst_mult_6_380 ;
wire Xd_0__inst_mult_7_372 ;
wire Xd_0__inst_mult_7_51_sumout ;
wire Xd_0__inst_mult_7_52 ;
wire Xd_0__inst_mult_7_53 ;
wire Xd_0__inst_mult_4_408 ;
wire Xd_0__inst_mult_5_372 ;
wire Xd_0__inst_mult_2_376 ;
wire Xd_0__inst_mult_3_372 ;
wire Xd_0__inst_mult_0_380 ;
wire Xd_0__inst_mult_0_55_sumout ;
wire Xd_0__inst_mult_0_56 ;
wire Xd_0__inst_mult_0_57 ;
wire Xd_0__inst_mult_1_380 ;
wire Xd_0__inst_mult_1_59_sumout ;
wire Xd_0__inst_mult_1_60 ;
wire Xd_0__inst_mult_1_61 ;
wire Xd_0__inst_mult_9_384 ;
wire Xd_0__inst_mult_9_385 ;
wire Xd_0__inst_mult_9_386 ;
wire Xd_0__inst_mult_9_388 ;
wire Xd_0__inst_mult_6_384 ;
wire Xd_0__inst_mult_6_385 ;
wire Xd_0__inst_mult_6_386 ;
wire Xd_0__inst_mult_6_388 ;
wire Xd_0__inst_mult_14_404 ;
wire Xd_0__inst_mult_14_405 ;
wire Xd_0__inst_mult_14_406 ;
wire Xd_0__inst_mult_14_408 ;
wire Xd_0__inst_mult_14_409 ;
wire Xd_0__inst_mult_14_410 ;
wire Xd_0__inst_mult_8_388 ;
wire Xd_0__inst_mult_8_389 ;
wire Xd_0__inst_mult_8_390 ;
wire Xd_0__inst_mult_8_392 ;
wire Xd_0__inst_mult_11_388 ;
wire Xd_0__inst_mult_11_389 ;
wire Xd_0__inst_mult_11_390 ;
wire Xd_0__inst_mult_11_392 ;
wire Xd_0__inst_mult_10_384 ;
wire Xd_0__inst_mult_10_385 ;
wire Xd_0__inst_mult_10_386 ;
wire Xd_0__inst_mult_10_388 ;
wire Xd_0__inst_mult_15_412 ;
wire Xd_0__inst_mult_15_413 ;
wire Xd_0__inst_mult_15_414 ;
wire Xd_0__inst_mult_13_388 ;
wire Xd_0__inst_mult_13_389 ;
wire Xd_0__inst_mult_13_390 ;
wire Xd_0__inst_mult_13_392 ;
wire Xd_0__inst_mult_15_416 ;
wire Xd_0__inst_mult_15_417 ;
wire Xd_0__inst_mult_15_418 ;
wire Xd_0__inst_mult_15_420 ;
wire Xd_0__inst_mult_12_408 ;
wire Xd_0__inst_mult_12_409 ;
wire Xd_0__inst_mult_12_410 ;
wire Xd_0__inst_mult_12_412 ;
wire Xd_0__inst_mult_12_416 ;
wire Xd_0__inst_mult_12_417 ;
wire Xd_0__inst_mult_12_418 ;
wire Xd_0__inst_mult_4_412 ;
wire Xd_0__inst_mult_4_413 ;
wire Xd_0__inst_mult_4_414 ;
wire Xd_0__inst_mult_12_420 ;
wire Xd_0__inst_mult_12_421 ;
wire Xd_0__inst_mult_12_422 ;
wire Xd_0__inst_mult_12_425 ;
wire Xd_0__inst_mult_12_426 ;
wire Xd_0__inst_mult_13_396 ;
wire Xd_0__inst_mult_13_397 ;
wire Xd_0__inst_mult_13_398 ;
wire Xd_0__inst_mult_13_401 ;
wire Xd_0__inst_mult_13_402 ;
wire Xd_0__inst_mult_14_412 ;
wire Xd_0__inst_mult_14_413 ;
wire Xd_0__inst_mult_14_414 ;
wire Xd_0__inst_mult_14_417 ;
wire Xd_0__inst_mult_14_418 ;
wire Xd_0__inst_mult_15_424 ;
wire Xd_0__inst_mult_15_425 ;
wire Xd_0__inst_mult_15_426 ;
wire Xd_0__inst_mult_15_429 ;
wire Xd_0__inst_mult_15_430 ;
wire Xd_0__inst_mult_10_392 ;
wire Xd_0__inst_mult_10_393 ;
wire Xd_0__inst_mult_10_394 ;
wire Xd_0__inst_mult_10_397 ;
wire Xd_0__inst_mult_10_398 ;
wire Xd_0__inst_mult_11_396 ;
wire Xd_0__inst_mult_11_397 ;
wire Xd_0__inst_mult_11_398 ;
wire Xd_0__inst_mult_11_401 ;
wire Xd_0__inst_mult_11_402 ;
wire Xd_0__inst_mult_8_396 ;
wire Xd_0__inst_mult_8_397 ;
wire Xd_0__inst_mult_8_398 ;
wire Xd_0__inst_mult_8_401 ;
wire Xd_0__inst_mult_8_402 ;
wire Xd_0__inst_mult_9_392 ;
wire Xd_0__inst_mult_9_393 ;
wire Xd_0__inst_mult_9_394 ;
wire Xd_0__inst_mult_9_397 ;
wire Xd_0__inst_mult_9_398 ;
wire Xd_0__inst_mult_6_392 ;
wire Xd_0__inst_mult_6_393 ;
wire Xd_0__inst_mult_6_394 ;
wire Xd_0__inst_mult_6_397 ;
wire Xd_0__inst_mult_6_398 ;
wire Xd_0__inst_mult_7_376 ;
wire Xd_0__inst_mult_7_377 ;
wire Xd_0__inst_mult_7_378 ;
wire Xd_0__inst_mult_7_380 ;
wire Xd_0__inst_mult_7_381 ;
wire Xd_0__inst_mult_7_382 ;
wire Xd_0__inst_mult_4_416 ;
wire Xd_0__inst_mult_4_417 ;
wire Xd_0__inst_mult_4_418 ;
wire Xd_0__inst_mult_4_420 ;
wire Xd_0__inst_mult_4_421 ;
wire Xd_0__inst_mult_4_422 ;
wire Xd_0__inst_mult_5_376 ;
wire Xd_0__inst_mult_5_377 ;
wire Xd_0__inst_mult_5_378 ;
wire Xd_0__inst_mult_5_380 ;
wire Xd_0__inst_mult_5_381 ;
wire Xd_0__inst_mult_5_382 ;
wire Xd_0__inst_mult_2_380 ;
wire Xd_0__inst_mult_2_381 ;
wire Xd_0__inst_mult_2_382 ;
wire Xd_0__inst_mult_2_384 ;
wire Xd_0__inst_mult_2_385 ;
wire Xd_0__inst_mult_2_386 ;
wire Xd_0__inst_mult_3_376 ;
wire Xd_0__inst_mult_3_377 ;
wire Xd_0__inst_mult_3_378 ;
wire Xd_0__inst_mult_3_380 ;
wire Xd_0__inst_mult_3_381 ;
wire Xd_0__inst_mult_3_382 ;
wire Xd_0__inst_mult_0_384 ;
wire Xd_0__inst_mult_0_385 ;
wire Xd_0__inst_mult_0_386 ;
wire Xd_0__inst_mult_1_384 ;
wire Xd_0__inst_mult_1_385 ;
wire Xd_0__inst_mult_1_386 ;
wire Xd_0__inst_mult_12_429 ;
wire Xd_0__inst_mult_12_430 ;
wire Xd_0__inst_mult_13_405 ;
wire Xd_0__inst_mult_13_406 ;
wire Xd_0__inst_mult_14_421 ;
wire Xd_0__inst_mult_14_422 ;
wire Xd_0__inst_mult_15_433 ;
wire Xd_0__inst_mult_15_434 ;
wire Xd_0__inst_mult_10_401 ;
wire Xd_0__inst_mult_10_402 ;
wire Xd_0__inst_mult_11_405 ;
wire Xd_0__inst_mult_11_406 ;
wire Xd_0__inst_mult_8_405 ;
wire Xd_0__inst_mult_8_406 ;
wire Xd_0__inst_mult_9_401 ;
wire Xd_0__inst_mult_9_402 ;
wire Xd_0__inst_mult_6_401 ;
wire Xd_0__inst_mult_6_402 ;
wire Xd_0__inst_mult_7_385 ;
wire Xd_0__inst_mult_7_386 ;
wire Xd_0__inst_mult_4_425 ;
wire Xd_0__inst_mult_4_426 ;
wire Xd_0__inst_mult_5_385 ;
wire Xd_0__inst_mult_5_386 ;
wire Xd_0__inst_mult_2_389 ;
wire Xd_0__inst_mult_2_390 ;
wire Xd_0__inst_mult_3_385 ;
wire Xd_0__inst_mult_3_386 ;
wire Xd_0__inst_mult_0_389 ;
wire Xd_0__inst_mult_0_390 ;
wire Xd_0__inst_mult_1_389 ;
wire Xd_0__inst_mult_1_390 ;
wire Xd_0__inst_mult_12_432 ;
wire Xd_0__inst_mult_12_433 ;
wire Xd_0__inst_mult_12_434 ;
wire Xd_0__inst_mult_12_436 ;
wire Xd_0__inst_mult_12_437 ;
wire Xd_0__inst_mult_12_438 ;
wire Xd_0__inst_mult_10_59_sumout ;
wire Xd_0__inst_mult_10_60 ;
wire Xd_0__inst_mult_10_61 ;
wire Xd_0__inst_mult_13_408 ;
wire Xd_0__inst_mult_13_409 ;
wire Xd_0__inst_mult_13_410 ;
wire Xd_0__inst_mult_13_412 ;
wire Xd_0__inst_mult_13_413 ;
wire Xd_0__inst_mult_13_414 ;
wire Xd_0__inst_mult_15_63_sumout ;
wire Xd_0__inst_mult_15_64 ;
wire Xd_0__inst_mult_15_65 ;
wire Xd_0__inst_mult_14_424 ;
wire Xd_0__inst_mult_14_425 ;
wire Xd_0__inst_mult_14_426 ;
wire Xd_0__inst_mult_14_428 ;
wire Xd_0__inst_mult_14_429 ;
wire Xd_0__inst_mult_14_430 ;
wire Xd_0__inst_mult_4_55_sumout ;
wire Xd_0__inst_mult_4_56 ;
wire Xd_0__inst_mult_4_57 ;
wire Xd_0__inst_mult_15_436 ;
wire Xd_0__inst_mult_15_437 ;
wire Xd_0__inst_mult_15_438 ;
wire Xd_0__inst_mult_15_440 ;
wire Xd_0__inst_mult_15_441 ;
wire Xd_0__inst_mult_15_442 ;
wire Xd_0__inst_mult_9_55_sumout ;
wire Xd_0__inst_mult_9_56 ;
wire Xd_0__inst_mult_9_57 ;
wire Xd_0__inst_mult_10_404 ;
wire Xd_0__inst_mult_10_405 ;
wire Xd_0__inst_mult_10_406 ;
wire Xd_0__inst_mult_10_408 ;
wire Xd_0__inst_mult_10_409 ;
wire Xd_0__inst_mult_10_410 ;
wire Xd_0__inst_mult_0_59_sumout ;
wire Xd_0__inst_mult_0_60 ;
wire Xd_0__inst_mult_0_61 ;
wire Xd_0__inst_mult_11_408 ;
wire Xd_0__inst_mult_11_409 ;
wire Xd_0__inst_mult_11_410 ;
wire Xd_0__inst_mult_11_412 ;
wire Xd_0__inst_mult_11_413 ;
wire Xd_0__inst_mult_11_414 ;
wire Xd_0__inst_mult_11_55_sumout ;
wire Xd_0__inst_mult_11_56 ;
wire Xd_0__inst_mult_11_57 ;
wire Xd_0__inst_mult_8_408 ;
wire Xd_0__inst_mult_8_409 ;
wire Xd_0__inst_mult_8_410 ;
wire Xd_0__inst_mult_8_412 ;
wire Xd_0__inst_mult_8_413 ;
wire Xd_0__inst_mult_8_414 ;
wire Xd_0__inst_mult_9_404 ;
wire Xd_0__inst_mult_9_405 ;
wire Xd_0__inst_mult_9_406 ;
wire Xd_0__inst_mult_9_408 ;
wire Xd_0__inst_mult_9_409 ;
wire Xd_0__inst_mult_9_410 ;
wire Xd_0__inst_mult_6_404 ;
wire Xd_0__inst_mult_6_405 ;
wire Xd_0__inst_mult_6_406 ;
wire Xd_0__inst_mult_6_408 ;
wire Xd_0__inst_mult_6_409 ;
wire Xd_0__inst_mult_6_410 ;
wire Xd_0__inst_mult_7_388 ;
wire Xd_0__inst_mult_7_389 ;
wire Xd_0__inst_mult_7_390 ;
wire Xd_0__inst_mult_7_392 ;
wire Xd_0__inst_mult_7_393 ;
wire Xd_0__inst_mult_7_394 ;
wire Xd_0__inst_mult_4_428 ;
wire Xd_0__inst_mult_4_429 ;
wire Xd_0__inst_mult_4_430 ;
wire Xd_0__inst_mult_4_432 ;
wire Xd_0__inst_mult_4_433 ;
wire Xd_0__inst_mult_4_434 ;
wire Xd_0__inst_mult_2_59_sumout ;
wire Xd_0__inst_mult_2_60 ;
wire Xd_0__inst_mult_2_61 ;
wire Xd_0__inst_mult_5_388 ;
wire Xd_0__inst_mult_5_389 ;
wire Xd_0__inst_mult_5_390 ;
wire Xd_0__inst_mult_5_392 ;
wire Xd_0__inst_mult_5_393 ;
wire Xd_0__inst_mult_5_394 ;
wire Xd_0__inst_mult_2_392 ;
wire Xd_0__inst_mult_2_393 ;
wire Xd_0__inst_mult_2_394 ;
wire Xd_0__inst_mult_2_396 ;
wire Xd_0__inst_mult_2_397 ;
wire Xd_0__inst_mult_2_398 ;
wire Xd_0__inst_mult_3_388 ;
wire Xd_0__inst_mult_3_389 ;
wire Xd_0__inst_mult_3_390 ;
wire Xd_0__inst_mult_3_392 ;
wire Xd_0__inst_mult_3_393 ;
wire Xd_0__inst_mult_3_394 ;
wire Xd_0__inst_mult_11_59_sumout ;
wire Xd_0__inst_mult_11_60 ;
wire Xd_0__inst_mult_11_61 ;
wire Xd_0__inst_mult_0_392 ;
wire Xd_0__inst_mult_0_393 ;
wire Xd_0__inst_mult_0_394 ;
wire Xd_0__inst_mult_0_396 ;
wire Xd_0__inst_mult_0_397 ;
wire Xd_0__inst_mult_0_398 ;
wire Xd_0__inst_mult_12_63_sumout ;
wire Xd_0__inst_mult_12_64 ;
wire Xd_0__inst_mult_12_65 ;
wire Xd_0__inst_mult_1_392 ;
wire Xd_0__inst_mult_1_393 ;
wire Xd_0__inst_mult_1_394 ;
wire Xd_0__inst_mult_1_396 ;
wire Xd_0__inst_mult_1_397 ;
wire Xd_0__inst_mult_1_398 ;
wire Xd_0__inst_mult_1_63_sumout ;
wire Xd_0__inst_mult_1_64 ;
wire Xd_0__inst_mult_1_65 ;
wire Xd_0__inst_mult_12_440 ;
wire Xd_0__inst_mult_12_441 ;
wire Xd_0__inst_mult_12_442 ;
wire Xd_0__inst_mult_12_444 ;
wire Xd_0__inst_mult_12_445 ;
wire Xd_0__inst_mult_12_446 ;
wire Xd_0__inst_mult_13_416 ;
wire Xd_0__inst_mult_13_417 ;
wire Xd_0__inst_mult_13_418 ;
wire Xd_0__inst_mult_13_420 ;
wire Xd_0__inst_mult_13_421 ;
wire Xd_0__inst_mult_13_422 ;
wire Xd_0__inst_mult_14_432 ;
wire Xd_0__inst_mult_14_433 ;
wire Xd_0__inst_mult_14_434 ;
wire Xd_0__inst_mult_14_436 ;
wire Xd_0__inst_mult_14_437 ;
wire Xd_0__inst_mult_14_438 ;
wire Xd_0__inst_mult_15_444 ;
wire Xd_0__inst_mult_15_445 ;
wire Xd_0__inst_mult_15_446 ;
wire Xd_0__inst_mult_15_448 ;
wire Xd_0__inst_mult_15_449 ;
wire Xd_0__inst_mult_15_450 ;
wire Xd_0__inst_mult_10_412 ;
wire Xd_0__inst_mult_10_413 ;
wire Xd_0__inst_mult_10_414 ;
wire Xd_0__inst_mult_10_416 ;
wire Xd_0__inst_mult_10_417 ;
wire Xd_0__inst_mult_10_418 ;
wire Xd_0__inst_mult_11_416 ;
wire Xd_0__inst_mult_11_417 ;
wire Xd_0__inst_mult_11_418 ;
wire Xd_0__inst_mult_11_420 ;
wire Xd_0__inst_mult_11_421 ;
wire Xd_0__inst_mult_11_422 ;
wire Xd_0__inst_mult_8_416 ;
wire Xd_0__inst_mult_8_417 ;
wire Xd_0__inst_mult_8_418 ;
wire Xd_0__inst_mult_8_420 ;
wire Xd_0__inst_mult_8_421 ;
wire Xd_0__inst_mult_8_422 ;
wire Xd_0__inst_mult_9_412 ;
wire Xd_0__inst_mult_9_413 ;
wire Xd_0__inst_mult_9_414 ;
wire Xd_0__inst_mult_9_416 ;
wire Xd_0__inst_mult_9_417 ;
wire Xd_0__inst_mult_9_418 ;
wire Xd_0__inst_mult_6_412 ;
wire Xd_0__inst_mult_6_413 ;
wire Xd_0__inst_mult_6_414 ;
wire Xd_0__inst_mult_6_416 ;
wire Xd_0__inst_mult_6_417 ;
wire Xd_0__inst_mult_6_418 ;
wire Xd_0__inst_mult_7_396 ;
wire Xd_0__inst_mult_7_397 ;
wire Xd_0__inst_mult_7_398 ;
wire Xd_0__inst_mult_7_400 ;
wire Xd_0__inst_mult_7_401 ;
wire Xd_0__inst_mult_7_402 ;
wire Xd_0__inst_mult_4_436 ;
wire Xd_0__inst_mult_4_437 ;
wire Xd_0__inst_mult_4_438 ;
wire Xd_0__inst_mult_4_440 ;
wire Xd_0__inst_mult_4_441 ;
wire Xd_0__inst_mult_4_442 ;
wire Xd_0__inst_mult_5_396 ;
wire Xd_0__inst_mult_5_397 ;
wire Xd_0__inst_mult_5_398 ;
wire Xd_0__inst_mult_5_400 ;
wire Xd_0__inst_mult_5_401 ;
wire Xd_0__inst_mult_5_402 ;
wire Xd_0__inst_mult_2_400 ;
wire Xd_0__inst_mult_2_401 ;
wire Xd_0__inst_mult_2_402 ;
wire Xd_0__inst_mult_2_404 ;
wire Xd_0__inst_mult_2_405 ;
wire Xd_0__inst_mult_2_406 ;
wire Xd_0__inst_mult_3_396 ;
wire Xd_0__inst_mult_3_397 ;
wire Xd_0__inst_mult_3_398 ;
wire Xd_0__inst_mult_3_400 ;
wire Xd_0__inst_mult_3_401 ;
wire Xd_0__inst_mult_3_402 ;
wire Xd_0__inst_mult_0_400 ;
wire Xd_0__inst_mult_0_401 ;
wire Xd_0__inst_mult_0_402 ;
wire Xd_0__inst_mult_0_404 ;
wire Xd_0__inst_mult_0_405 ;
wire Xd_0__inst_mult_0_406 ;
wire Xd_0__inst_mult_1_400 ;
wire Xd_0__inst_mult_1_401 ;
wire Xd_0__inst_mult_1_402 ;
wire Xd_0__inst_mult_1_404 ;
wire Xd_0__inst_mult_1_405 ;
wire Xd_0__inst_mult_1_406 ;
wire Xd_0__inst_mult_12_448 ;
wire Xd_0__inst_mult_12_449 ;
wire Xd_0__inst_mult_12_450 ;
wire Xd_0__inst_mult_12_452 ;
wire Xd_0__inst_mult_12_453 ;
wire Xd_0__inst_mult_12_454 ;
wire Xd_0__inst_mult_13_424 ;
wire Xd_0__inst_mult_13_425 ;
wire Xd_0__inst_mult_13_426 ;
wire Xd_0__inst_mult_13_428 ;
wire Xd_0__inst_mult_13_429 ;
wire Xd_0__inst_mult_13_430 ;
wire Xd_0__inst_mult_13_63_sumout ;
wire Xd_0__inst_mult_13_64 ;
wire Xd_0__inst_mult_13_65 ;
wire Xd_0__inst_mult_14_440 ;
wire Xd_0__inst_mult_14_441 ;
wire Xd_0__inst_mult_14_442 ;
wire Xd_0__inst_mult_14_444 ;
wire Xd_0__inst_mult_14_445 ;
wire Xd_0__inst_mult_14_446 ;
wire Xd_0__inst_mult_15_452 ;
wire Xd_0__inst_mult_15_453 ;
wire Xd_0__inst_mult_15_454 ;
wire Xd_0__inst_mult_15_456 ;
wire Xd_0__inst_mult_15_457 ;
wire Xd_0__inst_mult_15_458 ;
wire Xd_0__inst_mult_10_420 ;
wire Xd_0__inst_mult_10_421 ;
wire Xd_0__inst_mult_10_422 ;
wire Xd_0__inst_mult_10_424 ;
wire Xd_0__inst_mult_10_425 ;
wire Xd_0__inst_mult_10_426 ;
wire Xd_0__inst_mult_11_424 ;
wire Xd_0__inst_mult_11_425 ;
wire Xd_0__inst_mult_11_426 ;
wire Xd_0__inst_mult_11_428 ;
wire Xd_0__inst_mult_11_429 ;
wire Xd_0__inst_mult_11_430 ;
wire Xd_0__inst_mult_11_63_sumout ;
wire Xd_0__inst_mult_11_64 ;
wire Xd_0__inst_mult_11_65 ;
wire Xd_0__inst_mult_8_424 ;
wire Xd_0__inst_mult_8_425 ;
wire Xd_0__inst_mult_8_426 ;
wire Xd_0__inst_mult_8_428 ;
wire Xd_0__inst_mult_8_429 ;
wire Xd_0__inst_mult_8_430 ;
wire Xd_0__inst_mult_8_63_sumout ;
wire Xd_0__inst_mult_8_64 ;
wire Xd_0__inst_mult_8_65 ;
wire Xd_0__inst_mult_9_420 ;
wire Xd_0__inst_mult_9_421 ;
wire Xd_0__inst_mult_9_422 ;
wire Xd_0__inst_mult_9_424 ;
wire Xd_0__inst_mult_9_425 ;
wire Xd_0__inst_mult_9_426 ;
wire Xd_0__inst_mult_9_59_sumout ;
wire Xd_0__inst_mult_9_60 ;
wire Xd_0__inst_mult_9_61 ;
wire Xd_0__inst_mult_6_420 ;
wire Xd_0__inst_mult_6_421 ;
wire Xd_0__inst_mult_6_422 ;
wire Xd_0__inst_mult_6_424 ;
wire Xd_0__inst_mult_6_425 ;
wire Xd_0__inst_mult_6_426 ;
wire Xd_0__inst_mult_6_59_sumout ;
wire Xd_0__inst_mult_6_60 ;
wire Xd_0__inst_mult_6_61 ;
wire Xd_0__inst_mult_7_404 ;
wire Xd_0__inst_mult_7_405 ;
wire Xd_0__inst_mult_7_406 ;
wire Xd_0__inst_mult_7_408 ;
wire Xd_0__inst_mult_7_409 ;
wire Xd_0__inst_mult_7_410 ;
wire Xd_0__inst_mult_7_55_sumout ;
wire Xd_0__inst_mult_7_56 ;
wire Xd_0__inst_mult_7_57 ;
wire Xd_0__inst_mult_4_444 ;
wire Xd_0__inst_mult_4_445 ;
wire Xd_0__inst_mult_4_446 ;
wire Xd_0__inst_mult_4_448 ;
wire Xd_0__inst_mult_4_449 ;
wire Xd_0__inst_mult_4_450 ;
wire Xd_0__inst_mult_4_59_sumout ;
wire Xd_0__inst_mult_4_60 ;
wire Xd_0__inst_mult_4_61 ;
wire Xd_0__inst_mult_5_404 ;
wire Xd_0__inst_mult_5_405 ;
wire Xd_0__inst_mult_5_406 ;
wire Xd_0__inst_mult_5_408 ;
wire Xd_0__inst_mult_5_409 ;
wire Xd_0__inst_mult_5_410 ;
wire Xd_0__inst_mult_5_59_sumout ;
wire Xd_0__inst_mult_5_60 ;
wire Xd_0__inst_mult_5_61 ;
wire Xd_0__inst_mult_2_408 ;
wire Xd_0__inst_mult_2_409 ;
wire Xd_0__inst_mult_2_410 ;
wire Xd_0__inst_mult_2_412 ;
wire Xd_0__inst_mult_2_413 ;
wire Xd_0__inst_mult_2_414 ;
wire Xd_0__inst_mult_3_404 ;
wire Xd_0__inst_mult_3_405 ;
wire Xd_0__inst_mult_3_406 ;
wire Xd_0__inst_mult_3_408 ;
wire Xd_0__inst_mult_3_409 ;
wire Xd_0__inst_mult_3_410 ;
wire Xd_0__inst_mult_0_408 ;
wire Xd_0__inst_mult_0_409 ;
wire Xd_0__inst_mult_0_410 ;
wire Xd_0__inst_mult_0_412 ;
wire Xd_0__inst_mult_0_413 ;
wire Xd_0__inst_mult_0_414 ;
wire Xd_0__inst_mult_1_408 ;
wire Xd_0__inst_mult_1_409 ;
wire Xd_0__inst_mult_1_410 ;
wire Xd_0__inst_mult_1_412 ;
wire Xd_0__inst_mult_1_413 ;
wire Xd_0__inst_mult_1_414 ;
wire Xd_0__inst_mult_12_456 ;
wire Xd_0__inst_mult_12_457 ;
wire Xd_0__inst_mult_12_458 ;
wire Xd_0__inst_mult_12_460 ;
wire Xd_0__inst_mult_12_461 ;
wire Xd_0__inst_mult_12_462 ;
wire Xd_0__inst_mult_12_464 ;
wire Xd_0__inst_mult_12_465 ;
wire Xd_0__inst_mult_12_466 ;
wire Xd_0__inst_mult_12_469 ;
wire Xd_0__inst_mult_12_470 ;
wire Xd_0__inst_mult_13_432 ;
wire Xd_0__inst_mult_13_433 ;
wire Xd_0__inst_mult_13_434 ;
wire Xd_0__inst_mult_13_436 ;
wire Xd_0__inst_mult_13_437 ;
wire Xd_0__inst_mult_13_438 ;
wire Xd_0__inst_mult_13_440 ;
wire Xd_0__inst_mult_13_441 ;
wire Xd_0__inst_mult_13_442 ;
wire Xd_0__inst_mult_13_445 ;
wire Xd_0__inst_mult_13_446 ;
wire Xd_0__inst_mult_14_448 ;
wire Xd_0__inst_mult_14_449 ;
wire Xd_0__inst_mult_14_450 ;
wire Xd_0__inst_mult_14_452 ;
wire Xd_0__inst_mult_14_453 ;
wire Xd_0__inst_mult_14_454 ;
wire Xd_0__inst_mult_14_456 ;
wire Xd_0__inst_mult_14_457 ;
wire Xd_0__inst_mult_14_458 ;
wire Xd_0__inst_mult_14_461 ;
wire Xd_0__inst_mult_14_462 ;
wire Xd_0__inst_mult_15_460 ;
wire Xd_0__inst_mult_15_461 ;
wire Xd_0__inst_mult_15_462 ;
wire Xd_0__inst_mult_15_464 ;
wire Xd_0__inst_mult_15_465 ;
wire Xd_0__inst_mult_15_466 ;
wire Xd_0__inst_mult_15_468 ;
wire Xd_0__inst_mult_15_469 ;
wire Xd_0__inst_mult_15_470 ;
wire Xd_0__inst_mult_15_473 ;
wire Xd_0__inst_mult_15_474 ;
wire Xd_0__inst_mult_10_428 ;
wire Xd_0__inst_mult_10_429 ;
wire Xd_0__inst_mult_10_430 ;
wire Xd_0__inst_mult_10_432 ;
wire Xd_0__inst_mult_10_433 ;
wire Xd_0__inst_mult_10_434 ;
wire Xd_0__inst_mult_10_436 ;
wire Xd_0__inst_mult_10_437 ;
wire Xd_0__inst_mult_10_438 ;
wire Xd_0__inst_mult_10_441 ;
wire Xd_0__inst_mult_10_442 ;
wire Xd_0__inst_mult_11_432 ;
wire Xd_0__inst_mult_11_433 ;
wire Xd_0__inst_mult_11_434 ;
wire Xd_0__inst_mult_11_436 ;
wire Xd_0__inst_mult_11_437 ;
wire Xd_0__inst_mult_11_438 ;
wire Xd_0__inst_mult_11_440 ;
wire Xd_0__inst_mult_11_441 ;
wire Xd_0__inst_mult_11_442 ;
wire Xd_0__inst_mult_11_445 ;
wire Xd_0__inst_mult_11_446 ;
wire Xd_0__inst_mult_8_432 ;
wire Xd_0__inst_mult_8_433 ;
wire Xd_0__inst_mult_8_434 ;
wire Xd_0__inst_mult_8_436 ;
wire Xd_0__inst_mult_8_437 ;
wire Xd_0__inst_mult_8_438 ;
wire Xd_0__inst_mult_8_440 ;
wire Xd_0__inst_mult_8_441 ;
wire Xd_0__inst_mult_8_442 ;
wire Xd_0__inst_mult_8_445 ;
wire Xd_0__inst_mult_8_446 ;
wire Xd_0__inst_mult_9_428 ;
wire Xd_0__inst_mult_9_429 ;
wire Xd_0__inst_mult_9_430 ;
wire Xd_0__inst_mult_9_432 ;
wire Xd_0__inst_mult_9_433 ;
wire Xd_0__inst_mult_9_434 ;
wire Xd_0__inst_mult_9_63_sumout ;
wire Xd_0__inst_mult_9_64 ;
wire Xd_0__inst_mult_9_65 ;
wire Xd_0__inst_mult_9_436 ;
wire Xd_0__inst_mult_9_437 ;
wire Xd_0__inst_mult_9_438 ;
wire Xd_0__inst_mult_9_441 ;
wire Xd_0__inst_mult_9_442 ;
wire Xd_0__inst_mult_6_428 ;
wire Xd_0__inst_mult_6_429 ;
wire Xd_0__inst_mult_6_430 ;
wire Xd_0__inst_mult_6_432 ;
wire Xd_0__inst_mult_6_433 ;
wire Xd_0__inst_mult_6_434 ;
wire Xd_0__inst_mult_6_436 ;
wire Xd_0__inst_mult_6_437 ;
wire Xd_0__inst_mult_6_438 ;
wire Xd_0__inst_mult_6_441 ;
wire Xd_0__inst_mult_6_442 ;
wire Xd_0__inst_mult_7_412 ;
wire Xd_0__inst_mult_7_413 ;
wire Xd_0__inst_mult_7_414 ;
wire Xd_0__inst_mult_7_416 ;
wire Xd_0__inst_mult_7_417 ;
wire Xd_0__inst_mult_7_418 ;
wire Xd_0__inst_mult_7_59_sumout ;
wire Xd_0__inst_mult_7_60 ;
wire Xd_0__inst_mult_7_61 ;
wire Xd_0__inst_mult_7_420 ;
wire Xd_0__inst_mult_7_421 ;
wire Xd_0__inst_mult_7_422 ;
wire Xd_0__inst_mult_7_425 ;
wire Xd_0__inst_mult_7_426 ;
wire Xd_0__inst_mult_4_452 ;
wire Xd_0__inst_mult_4_453 ;
wire Xd_0__inst_mult_4_454 ;
wire Xd_0__inst_mult_4_456 ;
wire Xd_0__inst_mult_4_457 ;
wire Xd_0__inst_mult_4_458 ;
wire Xd_0__inst_mult_4_63_sumout ;
wire Xd_0__inst_mult_4_64 ;
wire Xd_0__inst_mult_4_65 ;
wire Xd_0__inst_mult_4_460 ;
wire Xd_0__inst_mult_4_461 ;
wire Xd_0__inst_mult_4_462 ;
wire Xd_0__inst_mult_4_465 ;
wire Xd_0__inst_mult_4_466 ;
wire Xd_0__inst_mult_5_412 ;
wire Xd_0__inst_mult_5_413 ;
wire Xd_0__inst_mult_5_414 ;
wire Xd_0__inst_mult_5_416 ;
wire Xd_0__inst_mult_5_417 ;
wire Xd_0__inst_mult_5_418 ;
wire Xd_0__inst_mult_5_63_sumout ;
wire Xd_0__inst_mult_5_64 ;
wire Xd_0__inst_mult_5_65 ;
wire Xd_0__inst_mult_5_420 ;
wire Xd_0__inst_mult_5_421 ;
wire Xd_0__inst_mult_5_422 ;
wire Xd_0__inst_mult_5_425 ;
wire Xd_0__inst_mult_5_426 ;
wire Xd_0__inst_mult_2_416 ;
wire Xd_0__inst_mult_2_417 ;
wire Xd_0__inst_mult_2_418 ;
wire Xd_0__inst_mult_2_420 ;
wire Xd_0__inst_mult_2_421 ;
wire Xd_0__inst_mult_2_422 ;
wire Xd_0__inst_mult_2_63_sumout ;
wire Xd_0__inst_mult_2_64 ;
wire Xd_0__inst_mult_2_65 ;
wire Xd_0__inst_mult_2_424 ;
wire Xd_0__inst_mult_2_425 ;
wire Xd_0__inst_mult_2_426 ;
wire Xd_0__inst_mult_2_429 ;
wire Xd_0__inst_mult_2_430 ;
wire Xd_0__inst_mult_3_412 ;
wire Xd_0__inst_mult_3_413 ;
wire Xd_0__inst_mult_3_414 ;
wire Xd_0__inst_mult_3_416 ;
wire Xd_0__inst_mult_3_417 ;
wire Xd_0__inst_mult_3_418 ;
wire Xd_0__inst_mult_3_420 ;
wire Xd_0__inst_mult_3_421 ;
wire Xd_0__inst_mult_3_422 ;
wire Xd_0__inst_mult_3_425 ;
wire Xd_0__inst_mult_3_426 ;
wire Xd_0__inst_mult_0_416 ;
wire Xd_0__inst_mult_0_417 ;
wire Xd_0__inst_mult_0_418 ;
wire Xd_0__inst_mult_0_420 ;
wire Xd_0__inst_mult_0_421 ;
wire Xd_0__inst_mult_0_422 ;
wire Xd_0__inst_mult_0_63_sumout ;
wire Xd_0__inst_mult_0_64 ;
wire Xd_0__inst_mult_0_65 ;
wire Xd_0__inst_mult_0_424 ;
wire Xd_0__inst_mult_0_425 ;
wire Xd_0__inst_mult_0_426 ;
wire Xd_0__inst_mult_0_429 ;
wire Xd_0__inst_mult_0_430 ;
wire Xd_0__inst_mult_1_416 ;
wire Xd_0__inst_mult_1_417 ;
wire Xd_0__inst_mult_1_418 ;
wire Xd_0__inst_mult_1_420 ;
wire Xd_0__inst_mult_1_421 ;
wire Xd_0__inst_mult_1_422 ;
wire Xd_0__inst_mult_1_67_sumout ;
wire Xd_0__inst_mult_1_68 ;
wire Xd_0__inst_mult_1_69 ;
wire Xd_0__inst_mult_1_424 ;
wire Xd_0__inst_mult_1_425 ;
wire Xd_0__inst_mult_1_426 ;
wire Xd_0__inst_mult_1_429 ;
wire Xd_0__inst_mult_1_430 ;
wire Xd_0__inst_mult_12_472 ;
wire Xd_0__inst_mult_12_473 ;
wire Xd_0__inst_mult_12_474 ;
wire Xd_0__inst_mult_12_476 ;
wire Xd_0__inst_mult_12_477 ;
wire Xd_0__inst_mult_12_478 ;
wire Xd_0__inst_mult_12_480 ;
wire Xd_0__inst_mult_12_481 ;
wire Xd_0__inst_mult_12_482 ;
wire Xd_0__inst_mult_12_484 ;
wire Xd_0__inst_mult_12_485 ;
wire Xd_0__inst_mult_12_486 ;
wire Xd_0__inst_mult_13_448 ;
wire Xd_0__inst_mult_13_449 ;
wire Xd_0__inst_mult_13_450 ;
wire Xd_0__inst_mult_13_452 ;
wire Xd_0__inst_mult_13_453 ;
wire Xd_0__inst_mult_13_454 ;
wire Xd_0__inst_mult_13_67_sumout ;
wire Xd_0__inst_mult_13_68 ;
wire Xd_0__inst_mult_13_69 ;
wire Xd_0__inst_mult_13_456 ;
wire Xd_0__inst_mult_13_457 ;
wire Xd_0__inst_mult_13_458 ;
wire Xd_0__inst_mult_13_460 ;
wire Xd_0__inst_mult_13_461 ;
wire Xd_0__inst_mult_13_462 ;
wire Xd_0__inst_mult_14_464 ;
wire Xd_0__inst_mult_14_465 ;
wire Xd_0__inst_mult_14_466 ;
wire Xd_0__inst_mult_14_468 ;
wire Xd_0__inst_mult_14_469 ;
wire Xd_0__inst_mult_14_470 ;
wire Xd_0__inst_mult_14_67_sumout ;
wire Xd_0__inst_mult_14_68 ;
wire Xd_0__inst_mult_14_69 ;
wire Xd_0__inst_mult_14_472 ;
wire Xd_0__inst_mult_14_473 ;
wire Xd_0__inst_mult_14_474 ;
wire Xd_0__inst_mult_14_476 ;
wire Xd_0__inst_mult_14_477 ;
wire Xd_0__inst_mult_14_478 ;
wire Xd_0__inst_mult_15_476 ;
wire Xd_0__inst_mult_15_477 ;
wire Xd_0__inst_mult_15_478 ;
wire Xd_0__inst_mult_15_480 ;
wire Xd_0__inst_mult_15_481 ;
wire Xd_0__inst_mult_15_482 ;
wire Xd_0__inst_mult_15_67_sumout ;
wire Xd_0__inst_mult_15_68 ;
wire Xd_0__inst_mult_15_69 ;
wire Xd_0__inst_mult_15_484 ;
wire Xd_0__inst_mult_15_485 ;
wire Xd_0__inst_mult_15_486 ;
wire Xd_0__inst_mult_15_488 ;
wire Xd_0__inst_mult_15_489 ;
wire Xd_0__inst_mult_15_490 ;
wire Xd_0__inst_mult_10_444 ;
wire Xd_0__inst_mult_10_445 ;
wire Xd_0__inst_mult_10_446 ;
wire Xd_0__inst_mult_10_448 ;
wire Xd_0__inst_mult_10_449 ;
wire Xd_0__inst_mult_10_450 ;
wire Xd_0__inst_mult_10_63_sumout ;
wire Xd_0__inst_mult_10_64 ;
wire Xd_0__inst_mult_10_65 ;
wire Xd_0__inst_mult_10_452 ;
wire Xd_0__inst_mult_10_453 ;
wire Xd_0__inst_mult_10_454 ;
wire Xd_0__inst_mult_10_456 ;
wire Xd_0__inst_mult_10_457 ;
wire Xd_0__inst_mult_10_458 ;
wire Xd_0__inst_mult_11_448 ;
wire Xd_0__inst_mult_11_449 ;
wire Xd_0__inst_mult_11_450 ;
wire Xd_0__inst_mult_11_452 ;
wire Xd_0__inst_mult_11_453 ;
wire Xd_0__inst_mult_11_454 ;
wire Xd_0__inst_mult_11_67_sumout ;
wire Xd_0__inst_mult_11_68 ;
wire Xd_0__inst_mult_11_69 ;
wire Xd_0__inst_mult_11_456 ;
wire Xd_0__inst_mult_11_457 ;
wire Xd_0__inst_mult_11_458 ;
wire Xd_0__inst_mult_11_460 ;
wire Xd_0__inst_mult_11_461 ;
wire Xd_0__inst_mult_11_462 ;
wire Xd_0__inst_mult_8_448 ;
wire Xd_0__inst_mult_8_449 ;
wire Xd_0__inst_mult_8_450 ;
wire Xd_0__inst_mult_8_452 ;
wire Xd_0__inst_mult_8_453 ;
wire Xd_0__inst_mult_8_454 ;
wire Xd_0__inst_mult_8_67_sumout ;
wire Xd_0__inst_mult_8_68 ;
wire Xd_0__inst_mult_8_69 ;
wire Xd_0__inst_mult_8_456 ;
wire Xd_0__inst_mult_8_457 ;
wire Xd_0__inst_mult_8_458 ;
wire Xd_0__inst_mult_8_460 ;
wire Xd_0__inst_mult_8_461 ;
wire Xd_0__inst_mult_8_462 ;
wire Xd_0__inst_mult_9_444 ;
wire Xd_0__inst_mult_9_445 ;
wire Xd_0__inst_mult_9_446 ;
wire Xd_0__inst_mult_9_448 ;
wire Xd_0__inst_mult_9_449 ;
wire Xd_0__inst_mult_9_450 ;
wire Xd_0__inst_mult_9_452 ;
wire Xd_0__inst_mult_9_453 ;
wire Xd_0__inst_mult_9_454 ;
wire Xd_0__inst_mult_9_456 ;
wire Xd_0__inst_mult_9_457 ;
wire Xd_0__inst_mult_9_458 ;
wire Xd_0__inst_mult_6_444 ;
wire Xd_0__inst_mult_6_445 ;
wire Xd_0__inst_mult_6_446 ;
wire Xd_0__inst_mult_6_448 ;
wire Xd_0__inst_mult_6_449 ;
wire Xd_0__inst_mult_6_450 ;
wire Xd_0__inst_mult_6_63_sumout ;
wire Xd_0__inst_mult_6_64 ;
wire Xd_0__inst_mult_6_65 ;
wire Xd_0__inst_mult_6_452 ;
wire Xd_0__inst_mult_6_453 ;
wire Xd_0__inst_mult_6_454 ;
wire Xd_0__inst_mult_6_456 ;
wire Xd_0__inst_mult_6_457 ;
wire Xd_0__inst_mult_6_458 ;
wire Xd_0__inst_mult_7_428 ;
wire Xd_0__inst_mult_7_429 ;
wire Xd_0__inst_mult_7_430 ;
wire Xd_0__inst_mult_7_432 ;
wire Xd_0__inst_mult_7_433 ;
wire Xd_0__inst_mult_7_434 ;
wire Xd_0__inst_mult_7_63_sumout ;
wire Xd_0__inst_mult_7_64 ;
wire Xd_0__inst_mult_7_65 ;
wire Xd_0__inst_mult_7_436 ;
wire Xd_0__inst_mult_7_437 ;
wire Xd_0__inst_mult_7_438 ;
wire Xd_0__inst_mult_7_440 ;
wire Xd_0__inst_mult_7_441 ;
wire Xd_0__inst_mult_7_442 ;
wire Xd_0__inst_mult_4_468 ;
wire Xd_0__inst_mult_4_469 ;
wire Xd_0__inst_mult_4_470 ;
wire Xd_0__inst_mult_4_472 ;
wire Xd_0__inst_mult_4_473 ;
wire Xd_0__inst_mult_4_474 ;
wire Xd_0__inst_mult_4_67_sumout ;
wire Xd_0__inst_mult_4_68 ;
wire Xd_0__inst_mult_4_69 ;
wire Xd_0__inst_mult_4_476 ;
wire Xd_0__inst_mult_4_477 ;
wire Xd_0__inst_mult_4_478 ;
wire Xd_0__inst_mult_4_480 ;
wire Xd_0__inst_mult_4_481 ;
wire Xd_0__inst_mult_4_482 ;
wire Xd_0__inst_mult_5_428 ;
wire Xd_0__inst_mult_5_429 ;
wire Xd_0__inst_mult_5_430 ;
wire Xd_0__inst_mult_5_432 ;
wire Xd_0__inst_mult_5_433 ;
wire Xd_0__inst_mult_5_434 ;
wire Xd_0__inst_mult_5_436 ;
wire Xd_0__inst_mult_5_437 ;
wire Xd_0__inst_mult_5_438 ;
wire Xd_0__inst_mult_5_440 ;
wire Xd_0__inst_mult_5_441 ;
wire Xd_0__inst_mult_5_442 ;
wire Xd_0__inst_mult_2_432 ;
wire Xd_0__inst_mult_2_433 ;
wire Xd_0__inst_mult_2_434 ;
wire Xd_0__inst_mult_2_436 ;
wire Xd_0__inst_mult_2_437 ;
wire Xd_0__inst_mult_2_438 ;
wire Xd_0__inst_mult_2_440 ;
wire Xd_0__inst_mult_2_441 ;
wire Xd_0__inst_mult_2_442 ;
wire Xd_0__inst_mult_2_444 ;
wire Xd_0__inst_mult_2_445 ;
wire Xd_0__inst_mult_2_446 ;
wire Xd_0__inst_mult_3_428 ;
wire Xd_0__inst_mult_3_429 ;
wire Xd_0__inst_mult_3_430 ;
wire Xd_0__inst_mult_3_432 ;
wire Xd_0__inst_mult_3_433 ;
wire Xd_0__inst_mult_3_434 ;
wire Xd_0__inst_mult_3_436 ;
wire Xd_0__inst_mult_3_437 ;
wire Xd_0__inst_mult_3_438 ;
wire Xd_0__inst_mult_3_440 ;
wire Xd_0__inst_mult_3_441 ;
wire Xd_0__inst_mult_3_442 ;
wire Xd_0__inst_mult_0_432 ;
wire Xd_0__inst_mult_0_433 ;
wire Xd_0__inst_mult_0_434 ;
wire Xd_0__inst_mult_0_436 ;
wire Xd_0__inst_mult_0_437 ;
wire Xd_0__inst_mult_0_438 ;
wire Xd_0__inst_mult_0_440 ;
wire Xd_0__inst_mult_0_441 ;
wire Xd_0__inst_mult_0_442 ;
wire Xd_0__inst_mult_0_444 ;
wire Xd_0__inst_mult_0_445 ;
wire Xd_0__inst_mult_0_446 ;
wire Xd_0__inst_mult_1_432 ;
wire Xd_0__inst_mult_1_433 ;
wire Xd_0__inst_mult_1_434 ;
wire Xd_0__inst_mult_1_436 ;
wire Xd_0__inst_mult_1_437 ;
wire Xd_0__inst_mult_1_438 ;
wire Xd_0__inst_mult_1_440 ;
wire Xd_0__inst_mult_1_441 ;
wire Xd_0__inst_mult_1_442 ;
wire Xd_0__inst_mult_1_444 ;
wire Xd_0__inst_mult_1_445 ;
wire Xd_0__inst_mult_1_446 ;
wire Xd_0__inst_mult_12_488 ;
wire Xd_0__inst_mult_12_489 ;
wire Xd_0__inst_mult_12_490 ;
wire Xd_0__inst_mult_12_492 ;
wire Xd_0__inst_mult_12_493 ;
wire Xd_0__inst_mult_12_494 ;
wire Xd_0__inst_mult_12_496 ;
wire Xd_0__inst_mult_12_497 ;
wire Xd_0__inst_mult_12_498 ;
wire Xd_0__inst_mult_12_500 ;
wire Xd_0__inst_mult_12_501 ;
wire Xd_0__inst_mult_12_502 ;
wire Xd_0__inst_mult_12_504 ;
wire Xd_0__inst_mult_12_505 ;
wire Xd_0__inst_mult_12_506 ;
wire Xd_0__inst_mult_13_464 ;
wire Xd_0__inst_mult_13_465 ;
wire Xd_0__inst_mult_13_466 ;
wire Xd_0__inst_mult_13_468 ;
wire Xd_0__inst_mult_13_469 ;
wire Xd_0__inst_mult_13_470 ;
wire Xd_0__inst_mult_13_472 ;
wire Xd_0__inst_mult_13_473 ;
wire Xd_0__inst_mult_13_474 ;
wire Xd_0__inst_mult_13_476 ;
wire Xd_0__inst_mult_13_477 ;
wire Xd_0__inst_mult_13_478 ;
wire Xd_0__inst_mult_13_480 ;
wire Xd_0__inst_mult_13_481 ;
wire Xd_0__inst_mult_13_482 ;
wire Xd_0__inst_mult_14_480 ;
wire Xd_0__inst_mult_14_481 ;
wire Xd_0__inst_mult_14_482 ;
wire Xd_0__inst_mult_14_484 ;
wire Xd_0__inst_mult_14_485 ;
wire Xd_0__inst_mult_14_486 ;
wire Xd_0__inst_mult_14_488 ;
wire Xd_0__inst_mult_14_489 ;
wire Xd_0__inst_mult_14_490 ;
wire Xd_0__inst_mult_15_492 ;
wire Xd_0__inst_mult_15_493 ;
wire Xd_0__inst_mult_15_494 ;
wire Xd_0__inst_mult_15_496 ;
wire Xd_0__inst_mult_15_497 ;
wire Xd_0__inst_mult_15_498 ;
wire Xd_0__inst_mult_15_500 ;
wire Xd_0__inst_mult_15_501 ;
wire Xd_0__inst_mult_15_502 ;
wire Xd_0__inst_mult_15_504 ;
wire Xd_0__inst_mult_15_505 ;
wire Xd_0__inst_mult_15_506 ;
wire Xd_0__inst_mult_15_508 ;
wire Xd_0__inst_mult_15_509 ;
wire Xd_0__inst_mult_15_510 ;
wire Xd_0__inst_mult_10_460 ;
wire Xd_0__inst_mult_10_461 ;
wire Xd_0__inst_mult_10_462 ;
wire Xd_0__inst_mult_10_464 ;
wire Xd_0__inst_mult_10_465 ;
wire Xd_0__inst_mult_10_466 ;
wire Xd_0__inst_mult_10_468 ;
wire Xd_0__inst_mult_10_469 ;
wire Xd_0__inst_mult_10_470 ;
wire Xd_0__inst_mult_10_472 ;
wire Xd_0__inst_mult_10_473 ;
wire Xd_0__inst_mult_10_474 ;
wire Xd_0__inst_mult_10_476 ;
wire Xd_0__inst_mult_10_477 ;
wire Xd_0__inst_mult_10_478 ;
wire Xd_0__inst_mult_11_464 ;
wire Xd_0__inst_mult_11_465 ;
wire Xd_0__inst_mult_11_466 ;
wire Xd_0__inst_mult_11_468 ;
wire Xd_0__inst_mult_11_469 ;
wire Xd_0__inst_mult_11_470 ;
wire Xd_0__inst_mult_11_472 ;
wire Xd_0__inst_mult_11_473 ;
wire Xd_0__inst_mult_11_474 ;
wire Xd_0__inst_mult_11_476 ;
wire Xd_0__inst_mult_11_477 ;
wire Xd_0__inst_mult_11_478 ;
wire Xd_0__inst_mult_11_480 ;
wire Xd_0__inst_mult_11_481 ;
wire Xd_0__inst_mult_11_482 ;
wire Xd_0__inst_mult_8_464 ;
wire Xd_0__inst_mult_8_465 ;
wire Xd_0__inst_mult_8_466 ;
wire Xd_0__inst_mult_8_468 ;
wire Xd_0__inst_mult_8_469 ;
wire Xd_0__inst_mult_8_470 ;
wire Xd_0__inst_mult_8_472 ;
wire Xd_0__inst_mult_8_473 ;
wire Xd_0__inst_mult_8_474 ;
wire Xd_0__inst_mult_8_476 ;
wire Xd_0__inst_mult_8_477 ;
wire Xd_0__inst_mult_8_478 ;
wire Xd_0__inst_mult_8_480 ;
wire Xd_0__inst_mult_8_481 ;
wire Xd_0__inst_mult_8_482 ;
wire Xd_0__inst_mult_9_460 ;
wire Xd_0__inst_mult_9_461 ;
wire Xd_0__inst_mult_9_462 ;
wire Xd_0__inst_mult_9_464 ;
wire Xd_0__inst_mult_9_465 ;
wire Xd_0__inst_mult_9_466 ;
wire Xd_0__inst_mult_9_468 ;
wire Xd_0__inst_mult_9_469 ;
wire Xd_0__inst_mult_9_470 ;
wire Xd_0__inst_mult_9_472 ;
wire Xd_0__inst_mult_9_473 ;
wire Xd_0__inst_mult_9_474 ;
wire Xd_0__inst_mult_9_476 ;
wire Xd_0__inst_mult_9_477 ;
wire Xd_0__inst_mult_9_478 ;
wire Xd_0__inst_mult_6_460 ;
wire Xd_0__inst_mult_6_461 ;
wire Xd_0__inst_mult_6_462 ;
wire Xd_0__inst_mult_6_464 ;
wire Xd_0__inst_mult_6_465 ;
wire Xd_0__inst_mult_6_466 ;
wire Xd_0__inst_mult_6_468 ;
wire Xd_0__inst_mult_6_469 ;
wire Xd_0__inst_mult_6_470 ;
wire Xd_0__inst_mult_6_472 ;
wire Xd_0__inst_mult_6_473 ;
wire Xd_0__inst_mult_6_474 ;
wire Xd_0__inst_mult_6_476 ;
wire Xd_0__inst_mult_6_477 ;
wire Xd_0__inst_mult_6_478 ;
wire Xd_0__inst_mult_7_444 ;
wire Xd_0__inst_mult_7_445 ;
wire Xd_0__inst_mult_7_446 ;
wire Xd_0__inst_mult_7_448 ;
wire Xd_0__inst_mult_7_449 ;
wire Xd_0__inst_mult_7_450 ;
wire Xd_0__inst_mult_7_452 ;
wire Xd_0__inst_mult_7_453 ;
wire Xd_0__inst_mult_7_454 ;
wire Xd_0__inst_mult_7_456 ;
wire Xd_0__inst_mult_7_457 ;
wire Xd_0__inst_mult_7_458 ;
wire Xd_0__inst_mult_7_460 ;
wire Xd_0__inst_mult_7_461 ;
wire Xd_0__inst_mult_7_462 ;
wire Xd_0__inst_mult_4_484 ;
wire Xd_0__inst_mult_4_485 ;
wire Xd_0__inst_mult_4_486 ;
wire Xd_0__inst_mult_4_488 ;
wire Xd_0__inst_mult_4_489 ;
wire Xd_0__inst_mult_4_490 ;
wire Xd_0__inst_mult_4_492 ;
wire Xd_0__inst_mult_4_493 ;
wire Xd_0__inst_mult_4_494 ;
wire Xd_0__inst_mult_4_496 ;
wire Xd_0__inst_mult_4_497 ;
wire Xd_0__inst_mult_4_498 ;
wire Xd_0__inst_mult_4_500 ;
wire Xd_0__inst_mult_4_501 ;
wire Xd_0__inst_mult_4_502 ;
wire Xd_0__inst_mult_5_444 ;
wire Xd_0__inst_mult_5_445 ;
wire Xd_0__inst_mult_5_446 ;
wire Xd_0__inst_mult_5_448 ;
wire Xd_0__inst_mult_5_449 ;
wire Xd_0__inst_mult_5_450 ;
wire Xd_0__inst_mult_5_452 ;
wire Xd_0__inst_mult_5_453 ;
wire Xd_0__inst_mult_5_454 ;
wire Xd_0__inst_mult_5_456 ;
wire Xd_0__inst_mult_5_457 ;
wire Xd_0__inst_mult_5_458 ;
wire Xd_0__inst_mult_5_460 ;
wire Xd_0__inst_mult_5_461 ;
wire Xd_0__inst_mult_5_462 ;
wire Xd_0__inst_mult_2_448 ;
wire Xd_0__inst_mult_2_449 ;
wire Xd_0__inst_mult_2_450 ;
wire Xd_0__inst_mult_2_452 ;
wire Xd_0__inst_mult_2_453 ;
wire Xd_0__inst_mult_2_454 ;
wire Xd_0__inst_mult_2_67_sumout ;
wire Xd_0__inst_mult_2_68 ;
wire Xd_0__inst_mult_2_69 ;
wire Xd_0__inst_mult_2_456 ;
wire Xd_0__inst_mult_2_457 ;
wire Xd_0__inst_mult_2_458 ;
wire Xd_0__inst_mult_2_460 ;
wire Xd_0__inst_mult_2_461 ;
wire Xd_0__inst_mult_2_462 ;
wire Xd_0__inst_mult_2_464 ;
wire Xd_0__inst_mult_2_465 ;
wire Xd_0__inst_mult_2_466 ;
wire Xd_0__inst_mult_3_444 ;
wire Xd_0__inst_mult_3_445 ;
wire Xd_0__inst_mult_3_446 ;
wire Xd_0__inst_mult_3_448 ;
wire Xd_0__inst_mult_3_449 ;
wire Xd_0__inst_mult_3_450 ;
wire Xd_0__inst_mult_3_63_sumout ;
wire Xd_0__inst_mult_3_64 ;
wire Xd_0__inst_mult_3_65 ;
wire Xd_0__inst_mult_3_452 ;
wire Xd_0__inst_mult_3_453 ;
wire Xd_0__inst_mult_3_454 ;
wire Xd_0__inst_mult_3_456 ;
wire Xd_0__inst_mult_3_457 ;
wire Xd_0__inst_mult_3_458 ;
wire Xd_0__inst_mult_3_460 ;
wire Xd_0__inst_mult_3_461 ;
wire Xd_0__inst_mult_3_462 ;
wire Xd_0__inst_mult_0_448 ;
wire Xd_0__inst_mult_0_449 ;
wire Xd_0__inst_mult_0_450 ;
wire Xd_0__inst_mult_0_452 ;
wire Xd_0__inst_mult_0_453 ;
wire Xd_0__inst_mult_0_454 ;
wire Xd_0__inst_mult_0_67_sumout ;
wire Xd_0__inst_mult_0_68 ;
wire Xd_0__inst_mult_0_69 ;
wire Xd_0__inst_mult_0_456 ;
wire Xd_0__inst_mult_0_457 ;
wire Xd_0__inst_mult_0_458 ;
wire Xd_0__inst_mult_0_460 ;
wire Xd_0__inst_mult_0_461 ;
wire Xd_0__inst_mult_0_462 ;
wire Xd_0__inst_mult_0_464 ;
wire Xd_0__inst_mult_0_465 ;
wire Xd_0__inst_mult_0_466 ;
wire Xd_0__inst_mult_1_448 ;
wire Xd_0__inst_mult_1_449 ;
wire Xd_0__inst_mult_1_450 ;
wire Xd_0__inst_mult_1_452 ;
wire Xd_0__inst_mult_1_453 ;
wire Xd_0__inst_mult_1_454 ;
wire Xd_0__inst_mult_1_456 ;
wire Xd_0__inst_mult_1_457 ;
wire Xd_0__inst_mult_1_458 ;
wire Xd_0__inst_mult_1_460 ;
wire Xd_0__inst_mult_1_461 ;
wire Xd_0__inst_mult_1_462 ;
wire Xd_0__inst_mult_1_464 ;
wire Xd_0__inst_mult_1_465 ;
wire Xd_0__inst_mult_1_466 ;
wire Xd_0__inst_mult_12_508 ;
wire Xd_0__inst_mult_12_509 ;
wire Xd_0__inst_mult_12_510 ;
wire Xd_0__inst_mult_12_512 ;
wire Xd_0__inst_mult_12_513 ;
wire Xd_0__inst_mult_12_514 ;
wire Xd_0__inst_mult_12_516 ;
wire Xd_0__inst_mult_12_517 ;
wire Xd_0__inst_mult_12_518 ;
wire Xd_0__inst_mult_12_520 ;
wire Xd_0__inst_mult_12_521 ;
wire Xd_0__inst_mult_12_522 ;
wire Xd_0__inst_mult_12_524 ;
wire Xd_0__inst_mult_12_525 ;
wire Xd_0__inst_mult_12_526 ;
wire Xd_0__inst_mult_13_484 ;
wire Xd_0__inst_mult_13_485 ;
wire Xd_0__inst_mult_13_486 ;
wire Xd_0__inst_mult_13_488 ;
wire Xd_0__inst_mult_13_489 ;
wire Xd_0__inst_mult_13_490 ;
wire Xd_0__inst_mult_13_492 ;
wire Xd_0__inst_mult_13_493 ;
wire Xd_0__inst_mult_13_494 ;
wire Xd_0__inst_mult_13_496 ;
wire Xd_0__inst_mult_13_497 ;
wire Xd_0__inst_mult_13_498 ;
wire Xd_0__inst_mult_13_500 ;
wire Xd_0__inst_mult_13_501 ;
wire Xd_0__inst_mult_13_502 ;
wire Xd_0__inst_mult_14_492 ;
wire Xd_0__inst_mult_14_493 ;
wire Xd_0__inst_mult_14_494 ;
wire Xd_0__inst_mult_14_496 ;
wire Xd_0__inst_mult_14_497 ;
wire Xd_0__inst_mult_14_498 ;
wire Xd_0__inst_mult_14_500 ;
wire Xd_0__inst_mult_14_501 ;
wire Xd_0__inst_mult_14_502 ;
wire Xd_0__inst_mult_15_512 ;
wire Xd_0__inst_mult_15_513 ;
wire Xd_0__inst_mult_15_514 ;
wire Xd_0__inst_mult_15_516 ;
wire Xd_0__inst_mult_15_517 ;
wire Xd_0__inst_mult_15_518 ;
wire Xd_0__inst_mult_15_520 ;
wire Xd_0__inst_mult_15_521 ;
wire Xd_0__inst_mult_15_522 ;
wire Xd_0__inst_mult_15_524 ;
wire Xd_0__inst_mult_15_525 ;
wire Xd_0__inst_mult_15_526 ;
wire Xd_0__inst_mult_15_528 ;
wire Xd_0__inst_mult_15_529 ;
wire Xd_0__inst_mult_15_530 ;
wire Xd_0__inst_mult_10_480 ;
wire Xd_0__inst_mult_10_481 ;
wire Xd_0__inst_mult_10_482 ;
wire Xd_0__inst_mult_10_484 ;
wire Xd_0__inst_mult_10_485 ;
wire Xd_0__inst_mult_10_486 ;
wire Xd_0__inst_mult_10_488 ;
wire Xd_0__inst_mult_10_489 ;
wire Xd_0__inst_mult_10_490 ;
wire Xd_0__inst_mult_10_492 ;
wire Xd_0__inst_mult_10_493 ;
wire Xd_0__inst_mult_10_494 ;
wire Xd_0__inst_mult_10_496 ;
wire Xd_0__inst_mult_10_497 ;
wire Xd_0__inst_mult_10_498 ;
wire Xd_0__inst_mult_11_484 ;
wire Xd_0__inst_mult_11_485 ;
wire Xd_0__inst_mult_11_486 ;
wire Xd_0__inst_mult_11_488 ;
wire Xd_0__inst_mult_11_489 ;
wire Xd_0__inst_mult_11_490 ;
wire Xd_0__inst_mult_11_492 ;
wire Xd_0__inst_mult_11_493 ;
wire Xd_0__inst_mult_11_494 ;
wire Xd_0__inst_mult_11_496 ;
wire Xd_0__inst_mult_11_497 ;
wire Xd_0__inst_mult_11_498 ;
wire Xd_0__inst_mult_11_500 ;
wire Xd_0__inst_mult_11_501 ;
wire Xd_0__inst_mult_11_502 ;
wire Xd_0__inst_mult_8_484 ;
wire Xd_0__inst_mult_8_485 ;
wire Xd_0__inst_mult_8_486 ;
wire Xd_0__inst_mult_8_488 ;
wire Xd_0__inst_mult_8_489 ;
wire Xd_0__inst_mult_8_490 ;
wire Xd_0__inst_mult_8_492 ;
wire Xd_0__inst_mult_8_493 ;
wire Xd_0__inst_mult_8_494 ;
wire Xd_0__inst_mult_8_496 ;
wire Xd_0__inst_mult_8_497 ;
wire Xd_0__inst_mult_8_498 ;
wire Xd_0__inst_mult_8_500 ;
wire Xd_0__inst_mult_8_501 ;
wire Xd_0__inst_mult_8_502 ;
wire Xd_0__inst_mult_9_480 ;
wire Xd_0__inst_mult_9_481 ;
wire Xd_0__inst_mult_9_482 ;
wire Xd_0__inst_mult_9_484 ;
wire Xd_0__inst_mult_9_485 ;
wire Xd_0__inst_mult_9_486 ;
wire Xd_0__inst_mult_9_488 ;
wire Xd_0__inst_mult_9_489 ;
wire Xd_0__inst_mult_9_490 ;
wire Xd_0__inst_mult_9_492 ;
wire Xd_0__inst_mult_9_493 ;
wire Xd_0__inst_mult_9_494 ;
wire Xd_0__inst_mult_9_496 ;
wire Xd_0__inst_mult_9_497 ;
wire Xd_0__inst_mult_9_498 ;
wire Xd_0__inst_mult_6_480 ;
wire Xd_0__inst_mult_6_481 ;
wire Xd_0__inst_mult_6_482 ;
wire Xd_0__inst_mult_6_484 ;
wire Xd_0__inst_mult_6_485 ;
wire Xd_0__inst_mult_6_486 ;
wire Xd_0__inst_mult_6_488 ;
wire Xd_0__inst_mult_6_489 ;
wire Xd_0__inst_mult_6_490 ;
wire Xd_0__inst_mult_6_492 ;
wire Xd_0__inst_mult_6_493 ;
wire Xd_0__inst_mult_6_494 ;
wire Xd_0__inst_mult_6_496 ;
wire Xd_0__inst_mult_6_497 ;
wire Xd_0__inst_mult_6_498 ;
wire Xd_0__inst_mult_7_464 ;
wire Xd_0__inst_mult_7_465 ;
wire Xd_0__inst_mult_7_466 ;
wire Xd_0__inst_mult_7_468 ;
wire Xd_0__inst_mult_7_469 ;
wire Xd_0__inst_mult_7_470 ;
wire Xd_0__inst_mult_7_472 ;
wire Xd_0__inst_mult_7_473 ;
wire Xd_0__inst_mult_7_474 ;
wire Xd_0__inst_mult_7_476 ;
wire Xd_0__inst_mult_7_477 ;
wire Xd_0__inst_mult_7_478 ;
wire Xd_0__inst_mult_7_480 ;
wire Xd_0__inst_mult_7_481 ;
wire Xd_0__inst_mult_7_482 ;
wire Xd_0__inst_mult_4_504 ;
wire Xd_0__inst_mult_4_505 ;
wire Xd_0__inst_mult_4_506 ;
wire Xd_0__inst_mult_4_508 ;
wire Xd_0__inst_mult_4_509 ;
wire Xd_0__inst_mult_4_510 ;
wire Xd_0__inst_mult_4_512 ;
wire Xd_0__inst_mult_4_513 ;
wire Xd_0__inst_mult_4_514 ;
wire Xd_0__inst_mult_4_516 ;
wire Xd_0__inst_mult_4_517 ;
wire Xd_0__inst_mult_4_518 ;
wire Xd_0__inst_mult_5_464 ;
wire Xd_0__inst_mult_5_465 ;
wire Xd_0__inst_mult_5_466 ;
wire Xd_0__inst_mult_5_468 ;
wire Xd_0__inst_mult_5_469 ;
wire Xd_0__inst_mult_5_470 ;
wire Xd_0__inst_mult_5_472 ;
wire Xd_0__inst_mult_5_473 ;
wire Xd_0__inst_mult_5_474 ;
wire Xd_0__inst_mult_5_476 ;
wire Xd_0__inst_mult_5_477 ;
wire Xd_0__inst_mult_5_478 ;
wire Xd_0__inst_mult_5_480 ;
wire Xd_0__inst_mult_5_481 ;
wire Xd_0__inst_mult_5_482 ;
wire Xd_0__inst_mult_2_468 ;
wire Xd_0__inst_mult_2_469 ;
wire Xd_0__inst_mult_2_470 ;
wire Xd_0__inst_mult_2_472 ;
wire Xd_0__inst_mult_2_473 ;
wire Xd_0__inst_mult_2_474 ;
wire Xd_0__inst_mult_2_476 ;
wire Xd_0__inst_mult_2_477 ;
wire Xd_0__inst_mult_2_478 ;
wire Xd_0__inst_mult_2_480 ;
wire Xd_0__inst_mult_2_481 ;
wire Xd_0__inst_mult_2_482 ;
wire Xd_0__inst_mult_2_484 ;
wire Xd_0__inst_mult_2_485 ;
wire Xd_0__inst_mult_2_486 ;
wire Xd_0__inst_mult_3_464 ;
wire Xd_0__inst_mult_3_465 ;
wire Xd_0__inst_mult_3_466 ;
wire Xd_0__inst_mult_3_468 ;
wire Xd_0__inst_mult_3_469 ;
wire Xd_0__inst_mult_3_470 ;
wire Xd_0__inst_mult_3_472 ;
wire Xd_0__inst_mult_3_473 ;
wire Xd_0__inst_mult_3_474 ;
wire Xd_0__inst_mult_3_476 ;
wire Xd_0__inst_mult_3_477 ;
wire Xd_0__inst_mult_3_478 ;
wire Xd_0__inst_mult_3_480 ;
wire Xd_0__inst_mult_3_481 ;
wire Xd_0__inst_mult_3_482 ;
wire Xd_0__inst_mult_0_468 ;
wire Xd_0__inst_mult_0_469 ;
wire Xd_0__inst_mult_0_470 ;
wire Xd_0__inst_mult_0_472 ;
wire Xd_0__inst_mult_0_473 ;
wire Xd_0__inst_mult_0_474 ;
wire Xd_0__inst_mult_0_476 ;
wire Xd_0__inst_mult_0_477 ;
wire Xd_0__inst_mult_0_478 ;
wire Xd_0__inst_mult_0_480 ;
wire Xd_0__inst_mult_0_481 ;
wire Xd_0__inst_mult_0_482 ;
wire Xd_0__inst_mult_0_484 ;
wire Xd_0__inst_mult_0_485 ;
wire Xd_0__inst_mult_0_486 ;
wire Xd_0__inst_mult_1_468 ;
wire Xd_0__inst_mult_1_469 ;
wire Xd_0__inst_mult_1_470 ;
wire Xd_0__inst_mult_1_472 ;
wire Xd_0__inst_mult_1_473 ;
wire Xd_0__inst_mult_1_474 ;
wire Xd_0__inst_mult_1_476 ;
wire Xd_0__inst_mult_1_477 ;
wire Xd_0__inst_mult_1_478 ;
wire Xd_0__inst_mult_1_480 ;
wire Xd_0__inst_mult_1_481 ;
wire Xd_0__inst_mult_1_482 ;
wire Xd_0__inst_mult_1_484 ;
wire Xd_0__inst_mult_1_485 ;
wire Xd_0__inst_mult_1_486 ;
wire Xd_0__inst_mult_12_528 ;
wire Xd_0__inst_mult_12_529 ;
wire Xd_0__inst_mult_12_530 ;
wire Xd_0__inst_mult_12_532 ;
wire Xd_0__inst_mult_12_533 ;
wire Xd_0__inst_mult_12_534 ;
wire Xd_0__inst_mult_12_536 ;
wire Xd_0__inst_mult_12_537 ;
wire Xd_0__inst_mult_12_538 ;
wire Xd_0__inst_mult_13_504 ;
wire Xd_0__inst_mult_13_505 ;
wire Xd_0__inst_mult_13_506 ;
wire Xd_0__inst_mult_13_508 ;
wire Xd_0__inst_mult_13_509 ;
wire Xd_0__inst_mult_13_510 ;
wire Xd_0__inst_mult_13_512 ;
wire Xd_0__inst_mult_13_513 ;
wire Xd_0__inst_mult_13_514 ;
wire Xd_0__inst_mult_14_504 ;
wire Xd_0__inst_mult_14_505 ;
wire Xd_0__inst_mult_14_506 ;
wire Xd_0__inst_mult_14_508 ;
wire Xd_0__inst_mult_14_509 ;
wire Xd_0__inst_mult_14_510 ;
wire Xd_0__inst_mult_14_512 ;
wire Xd_0__inst_mult_14_513 ;
wire Xd_0__inst_mult_14_514 ;
wire Xd_0__inst_mult_15_532 ;
wire Xd_0__inst_mult_15_533 ;
wire Xd_0__inst_mult_15_534 ;
wire Xd_0__inst_mult_15_536 ;
wire Xd_0__inst_mult_15_537 ;
wire Xd_0__inst_mult_15_538 ;
wire Xd_0__inst_mult_15_540 ;
wire Xd_0__inst_mult_15_541 ;
wire Xd_0__inst_mult_15_542 ;
wire Xd_0__inst_mult_10_500 ;
wire Xd_0__inst_mult_10_501 ;
wire Xd_0__inst_mult_10_502 ;
wire Xd_0__inst_mult_10_504 ;
wire Xd_0__inst_mult_10_505 ;
wire Xd_0__inst_mult_10_506 ;
wire Xd_0__inst_mult_10_508 ;
wire Xd_0__inst_mult_10_509 ;
wire Xd_0__inst_mult_10_510 ;
wire Xd_0__inst_mult_11_504 ;
wire Xd_0__inst_mult_11_505 ;
wire Xd_0__inst_mult_11_506 ;
wire Xd_0__inst_mult_11_508 ;
wire Xd_0__inst_mult_11_509 ;
wire Xd_0__inst_mult_11_510 ;
wire Xd_0__inst_mult_11_512 ;
wire Xd_0__inst_mult_11_513 ;
wire Xd_0__inst_mult_11_514 ;
wire Xd_0__inst_mult_8_504 ;
wire Xd_0__inst_mult_8_505 ;
wire Xd_0__inst_mult_8_506 ;
wire Xd_0__inst_mult_8_508 ;
wire Xd_0__inst_mult_8_509 ;
wire Xd_0__inst_mult_8_510 ;
wire Xd_0__inst_mult_8_512 ;
wire Xd_0__inst_mult_8_513 ;
wire Xd_0__inst_mult_8_514 ;
wire Xd_0__inst_mult_9_500 ;
wire Xd_0__inst_mult_9_501 ;
wire Xd_0__inst_mult_9_502 ;
wire Xd_0__inst_mult_9_504 ;
wire Xd_0__inst_mult_9_505 ;
wire Xd_0__inst_mult_9_506 ;
wire Xd_0__inst_mult_9_508 ;
wire Xd_0__inst_mult_9_509 ;
wire Xd_0__inst_mult_9_510 ;
wire Xd_0__inst_mult_6_500 ;
wire Xd_0__inst_mult_6_501 ;
wire Xd_0__inst_mult_6_502 ;
wire Xd_0__inst_mult_6_504 ;
wire Xd_0__inst_mult_6_505 ;
wire Xd_0__inst_mult_6_506 ;
wire Xd_0__inst_mult_6_508 ;
wire Xd_0__inst_mult_6_509 ;
wire Xd_0__inst_mult_6_510 ;
wire Xd_0__inst_mult_7_484 ;
wire Xd_0__inst_mult_7_488 ;
wire Xd_0__inst_mult_7_489 ;
wire Xd_0__inst_mult_7_490 ;
wire Xd_0__inst_mult_7_492 ;
wire Xd_0__inst_mult_7_493 ;
wire Xd_0__inst_mult_7_494 ;
wire Xd_0__inst_mult_7_496 ;
wire Xd_0__inst_mult_7_497 ;
wire Xd_0__inst_mult_7_498 ;
wire Xd_0__inst_mult_7_500 ;
wire Xd_0__inst_mult_7_501 ;
wire Xd_0__inst_mult_7_502 ;
wire Xd_0__inst_mult_4_520 ;
wire Xd_0__inst_mult_4_524 ;
wire Xd_0__inst_mult_4_525 ;
wire Xd_0__inst_mult_4_526 ;
wire Xd_0__inst_mult_4_528 ;
wire Xd_0__inst_mult_4_529 ;
wire Xd_0__inst_mult_4_530 ;
wire Xd_0__inst_mult_4_532 ;
wire Xd_0__inst_mult_4_533 ;
wire Xd_0__inst_mult_4_534 ;
wire Xd_0__inst_mult_5_484 ;
wire Xd_0__inst_mult_5_488 ;
wire Xd_0__inst_mult_5_489 ;
wire Xd_0__inst_mult_5_490 ;
wire Xd_0__inst_mult_5_492 ;
wire Xd_0__inst_mult_5_493 ;
wire Xd_0__inst_mult_5_494 ;
wire Xd_0__inst_mult_5_496 ;
wire Xd_0__inst_mult_5_497 ;
wire Xd_0__inst_mult_5_498 ;
wire Xd_0__inst_mult_5_500 ;
wire Xd_0__inst_mult_5_501 ;
wire Xd_0__inst_mult_5_502 ;
wire Xd_0__inst_mult_2_488 ;
wire Xd_0__inst_mult_2_492 ;
wire Xd_0__inst_mult_2_493 ;
wire Xd_0__inst_mult_2_494 ;
wire Xd_0__inst_mult_2_496 ;
wire Xd_0__inst_mult_2_497 ;
wire Xd_0__inst_mult_2_498 ;
wire Xd_0__inst_mult_2_500 ;
wire Xd_0__inst_mult_2_501 ;
wire Xd_0__inst_mult_2_502 ;
wire Xd_0__inst_mult_2_504 ;
wire Xd_0__inst_mult_2_505 ;
wire Xd_0__inst_mult_2_506 ;
wire Xd_0__inst_mult_3_484 ;
wire Xd_0__inst_mult_3_488 ;
wire Xd_0__inst_mult_3_489 ;
wire Xd_0__inst_mult_3_490 ;
wire Xd_0__inst_mult_3_492 ;
wire Xd_0__inst_mult_3_493 ;
wire Xd_0__inst_mult_3_494 ;
wire Xd_0__inst_mult_3_496 ;
wire Xd_0__inst_mult_3_497 ;
wire Xd_0__inst_mult_3_498 ;
wire Xd_0__inst_mult_3_500 ;
wire Xd_0__inst_mult_3_501 ;
wire Xd_0__inst_mult_3_502 ;
wire Xd_0__inst_mult_0_488 ;
wire Xd_0__inst_mult_0_492 ;
wire Xd_0__inst_mult_0_493 ;
wire Xd_0__inst_mult_0_494 ;
wire Xd_0__inst_mult_0_496 ;
wire Xd_0__inst_mult_0_497 ;
wire Xd_0__inst_mult_0_498 ;
wire Xd_0__inst_mult_0_500 ;
wire Xd_0__inst_mult_0_501 ;
wire Xd_0__inst_mult_0_502 ;
wire Xd_0__inst_mult_0_504 ;
wire Xd_0__inst_mult_0_505 ;
wire Xd_0__inst_mult_0_506 ;
wire Xd_0__inst_mult_1_488 ;
wire Xd_0__inst_mult_1_492 ;
wire Xd_0__inst_mult_1_493 ;
wire Xd_0__inst_mult_1_494 ;
wire Xd_0__inst_mult_1_496 ;
wire Xd_0__inst_mult_1_497 ;
wire Xd_0__inst_mult_1_498 ;
wire Xd_0__inst_mult_1_500 ;
wire Xd_0__inst_mult_1_501 ;
wire Xd_0__inst_mult_1_502 ;
wire Xd_0__inst_mult_1_504 ;
wire Xd_0__inst_mult_1_505 ;
wire Xd_0__inst_mult_1_506 ;
wire Xd_0__inst_mult_12_540 ;
wire Xd_0__inst_mult_12_541 ;
wire Xd_0__inst_mult_12_542 ;
wire Xd_0__inst_mult_12_544 ;
wire Xd_0__inst_mult_12_545 ;
wire Xd_0__inst_mult_12_546 ;
wire Xd_0__inst_mult_13_516 ;
wire Xd_0__inst_mult_13_517 ;
wire Xd_0__inst_mult_13_518 ;
wire Xd_0__inst_mult_13_520 ;
wire Xd_0__inst_mult_13_521 ;
wire Xd_0__inst_mult_13_522 ;
wire Xd_0__inst_mult_13_524 ;
wire Xd_0__inst_mult_13_525 ;
wire Xd_0__inst_mult_13_526 ;
wire Xd_0__inst_mult_14_516 ;
wire Xd_0__inst_mult_14_517 ;
wire Xd_0__inst_mult_14_518 ;
wire Xd_0__inst_mult_14_520 ;
wire Xd_0__inst_mult_14_521 ;
wire Xd_0__inst_mult_14_522 ;
wire Xd_0__inst_mult_14_524 ;
wire Xd_0__inst_mult_14_525 ;
wire Xd_0__inst_mult_14_526 ;
wire Xd_0__inst_mult_15_544 ;
wire Xd_0__inst_mult_15_545 ;
wire Xd_0__inst_mult_15_546 ;
wire Xd_0__inst_mult_15_548 ;
wire Xd_0__inst_mult_15_549 ;
wire Xd_0__inst_mult_15_550 ;
wire Xd_0__inst_mult_10_512 ;
wire Xd_0__inst_mult_10_513 ;
wire Xd_0__inst_mult_10_514 ;
wire Xd_0__inst_mult_10_516 ;
wire Xd_0__inst_mult_10_517 ;
wire Xd_0__inst_mult_10_518 ;
wire Xd_0__inst_mult_10_520 ;
wire Xd_0__inst_mult_10_521 ;
wire Xd_0__inst_mult_10_522 ;
wire Xd_0__inst_mult_11_516 ;
wire Xd_0__inst_mult_11_517 ;
wire Xd_0__inst_mult_11_518 ;
wire Xd_0__inst_mult_11_520 ;
wire Xd_0__inst_mult_11_521 ;
wire Xd_0__inst_mult_11_522 ;
wire Xd_0__inst_mult_11_524 ;
wire Xd_0__inst_mult_11_525 ;
wire Xd_0__inst_mult_11_526 ;
wire Xd_0__inst_mult_8_516 ;
wire Xd_0__inst_mult_8_517 ;
wire Xd_0__inst_mult_8_518 ;
wire Xd_0__inst_mult_8_520 ;
wire Xd_0__inst_mult_8_521 ;
wire Xd_0__inst_mult_8_522 ;
wire Xd_0__inst_mult_8_524 ;
wire Xd_0__inst_mult_8_525 ;
wire Xd_0__inst_mult_8_526 ;
wire Xd_0__inst_mult_9_512 ;
wire Xd_0__inst_mult_9_513 ;
wire Xd_0__inst_mult_9_514 ;
wire Xd_0__inst_mult_9_516 ;
wire Xd_0__inst_mult_9_517 ;
wire Xd_0__inst_mult_9_518 ;
wire Xd_0__inst_mult_9_520 ;
wire Xd_0__inst_mult_9_521 ;
wire Xd_0__inst_mult_9_522 ;
wire Xd_0__inst_mult_6_512 ;
wire Xd_0__inst_mult_6_513 ;
wire Xd_0__inst_mult_6_514 ;
wire Xd_0__inst_mult_6_516 ;
wire Xd_0__inst_mult_6_517 ;
wire Xd_0__inst_mult_6_518 ;
wire Xd_0__inst_mult_6_520 ;
wire Xd_0__inst_mult_6_521 ;
wire Xd_0__inst_mult_6_522 ;
wire Xd_0__inst_mult_7_504 ;
wire Xd_0__inst_mult_7_505 ;
wire Xd_0__inst_mult_7_506 ;
wire Xd_0__inst_mult_7_508 ;
wire Xd_0__inst_mult_7_509 ;
wire Xd_0__inst_mult_7_510 ;
wire Xd_0__inst_mult_7_512 ;
wire Xd_0__inst_mult_7_513 ;
wire Xd_0__inst_mult_7_514 ;
wire Xd_0__inst_mult_7_516 ;
wire Xd_0__inst_mult_7_517 ;
wire Xd_0__inst_mult_7_518 ;
wire Xd_0__inst_mult_4_536 ;
wire Xd_0__inst_mult_4_537 ;
wire Xd_0__inst_mult_4_538 ;
wire Xd_0__inst_mult_4_540 ;
wire Xd_0__inst_mult_4_541 ;
wire Xd_0__inst_mult_4_542 ;
wire Xd_0__inst_mult_4_544 ;
wire Xd_0__inst_mult_4_545 ;
wire Xd_0__inst_mult_4_546 ;
wire Xd_0__inst_mult_5_504 ;
wire Xd_0__inst_mult_5_505 ;
wire Xd_0__inst_mult_5_506 ;
wire Xd_0__inst_mult_5_508 ;
wire Xd_0__inst_mult_5_509 ;
wire Xd_0__inst_mult_5_510 ;
wire Xd_0__inst_mult_5_512 ;
wire Xd_0__inst_mult_5_513 ;
wire Xd_0__inst_mult_5_514 ;
wire Xd_0__inst_mult_5_516 ;
wire Xd_0__inst_mult_5_517 ;
wire Xd_0__inst_mult_5_518 ;
wire Xd_0__inst_mult_2_508 ;
wire Xd_0__inst_mult_2_509 ;
wire Xd_0__inst_mult_2_510 ;
wire Xd_0__inst_mult_2_512 ;
wire Xd_0__inst_mult_2_513 ;
wire Xd_0__inst_mult_2_514 ;
wire Xd_0__inst_mult_2_516 ;
wire Xd_0__inst_mult_2_517 ;
wire Xd_0__inst_mult_2_518 ;
wire Xd_0__inst_mult_2_520 ;
wire Xd_0__inst_mult_2_521 ;
wire Xd_0__inst_mult_2_522 ;
wire Xd_0__inst_mult_3_504 ;
wire Xd_0__inst_mult_3_505 ;
wire Xd_0__inst_mult_3_506 ;
wire Xd_0__inst_mult_3_508 ;
wire Xd_0__inst_mult_3_509 ;
wire Xd_0__inst_mult_3_510 ;
wire Xd_0__inst_mult_3_512 ;
wire Xd_0__inst_mult_3_513 ;
wire Xd_0__inst_mult_3_514 ;
wire Xd_0__inst_mult_3_516 ;
wire Xd_0__inst_mult_3_517 ;
wire Xd_0__inst_mult_3_518 ;
wire Xd_0__inst_mult_0_508 ;
wire Xd_0__inst_mult_0_509 ;
wire Xd_0__inst_mult_0_510 ;
wire Xd_0__inst_mult_0_512 ;
wire Xd_0__inst_mult_0_513 ;
wire Xd_0__inst_mult_0_514 ;
wire Xd_0__inst_mult_0_516 ;
wire Xd_0__inst_mult_0_517 ;
wire Xd_0__inst_mult_0_518 ;
wire Xd_0__inst_mult_0_520 ;
wire Xd_0__inst_mult_0_521 ;
wire Xd_0__inst_mult_0_522 ;
wire Xd_0__inst_mult_1_508 ;
wire Xd_0__inst_mult_1_509 ;
wire Xd_0__inst_mult_1_510 ;
wire Xd_0__inst_mult_1_512 ;
wire Xd_0__inst_mult_1_513 ;
wire Xd_0__inst_mult_1_514 ;
wire Xd_0__inst_mult_1_516 ;
wire Xd_0__inst_mult_1_517 ;
wire Xd_0__inst_mult_1_518 ;
wire Xd_0__inst_mult_1_520 ;
wire Xd_0__inst_mult_1_521 ;
wire Xd_0__inst_mult_1_522 ;
wire Xd_0__inst_mult_12_548 ;
wire Xd_0__inst_mult_12_549 ;
wire Xd_0__inst_mult_12_550 ;
wire Xd_0__inst_mult_12_552 ;
wire Xd_0__inst_mult_12_553 ;
wire Xd_0__inst_mult_12_554 ;
wire Xd_0__inst_mult_13_528 ;
wire Xd_0__inst_mult_13_529 ;
wire Xd_0__inst_mult_13_530 ;
wire Xd_0__inst_mult_13_532 ;
wire Xd_0__inst_mult_13_533 ;
wire Xd_0__inst_mult_13_534 ;
wire Xd_0__inst_mult_13_536 ;
wire Xd_0__inst_mult_13_537 ;
wire Xd_0__inst_mult_13_538 ;
wire Xd_0__inst_mult_14_528 ;
wire Xd_0__inst_mult_14_529 ;
wire Xd_0__inst_mult_14_530 ;
wire Xd_0__inst_mult_14_532 ;
wire Xd_0__inst_mult_14_533 ;
wire Xd_0__inst_mult_14_534 ;
wire Xd_0__inst_mult_14_536 ;
wire Xd_0__inst_mult_14_537 ;
wire Xd_0__inst_mult_14_538 ;
wire Xd_0__inst_mult_15_552 ;
wire Xd_0__inst_mult_15_553 ;
wire Xd_0__inst_mult_15_554 ;
wire Xd_0__inst_mult_15_556 ;
wire Xd_0__inst_mult_15_557 ;
wire Xd_0__inst_mult_15_558 ;
wire Xd_0__inst_mult_10_524 ;
wire Xd_0__inst_mult_10_525 ;
wire Xd_0__inst_mult_10_526 ;
wire Xd_0__inst_mult_10_528 ;
wire Xd_0__inst_mult_10_529 ;
wire Xd_0__inst_mult_10_530 ;
wire Xd_0__inst_mult_10_532 ;
wire Xd_0__inst_mult_10_533 ;
wire Xd_0__inst_mult_10_534 ;
wire Xd_0__inst_mult_11_528 ;
wire Xd_0__inst_mult_11_529 ;
wire Xd_0__inst_mult_11_530 ;
wire Xd_0__inst_mult_11_532 ;
wire Xd_0__inst_mult_11_533 ;
wire Xd_0__inst_mult_11_534 ;
wire Xd_0__inst_mult_11_536 ;
wire Xd_0__inst_mult_11_537 ;
wire Xd_0__inst_mult_11_538 ;
wire Xd_0__inst_mult_8_528 ;
wire Xd_0__inst_mult_8_529 ;
wire Xd_0__inst_mult_8_530 ;
wire Xd_0__inst_mult_8_532 ;
wire Xd_0__inst_mult_8_533 ;
wire Xd_0__inst_mult_8_534 ;
wire Xd_0__inst_mult_8_536 ;
wire Xd_0__inst_mult_8_537 ;
wire Xd_0__inst_mult_8_538 ;
wire Xd_0__inst_mult_9_524 ;
wire Xd_0__inst_mult_9_525 ;
wire Xd_0__inst_mult_9_526 ;
wire Xd_0__inst_mult_9_528 ;
wire Xd_0__inst_mult_9_529 ;
wire Xd_0__inst_mult_9_530 ;
wire Xd_0__inst_mult_9_532 ;
wire Xd_0__inst_mult_9_533 ;
wire Xd_0__inst_mult_9_534 ;
wire Xd_0__inst_mult_6_524 ;
wire Xd_0__inst_mult_6_525 ;
wire Xd_0__inst_mult_6_526 ;
wire Xd_0__inst_mult_6_528 ;
wire Xd_0__inst_mult_6_529 ;
wire Xd_0__inst_mult_6_530 ;
wire Xd_0__inst_mult_6_532 ;
wire Xd_0__inst_mult_6_533 ;
wire Xd_0__inst_mult_6_534 ;
wire Xd_0__inst_mult_7_520 ;
wire Xd_0__inst_mult_7_524 ;
wire Xd_0__inst_mult_7_525 ;
wire Xd_0__inst_mult_7_526 ;
wire Xd_0__inst_mult_7_528 ;
wire Xd_0__inst_mult_7_529 ;
wire Xd_0__inst_mult_7_530 ;
wire Xd_0__inst_mult_7_532 ;
wire Xd_0__inst_mult_7_533 ;
wire Xd_0__inst_mult_7_534 ;
wire Xd_0__inst_mult_4_548 ;
wire Xd_0__inst_mult_4_552 ;
wire Xd_0__inst_mult_4_553 ;
wire Xd_0__inst_mult_4_554 ;
wire Xd_0__inst_mult_4_556 ;
wire Xd_0__inst_mult_4_557 ;
wire Xd_0__inst_mult_4_558 ;
wire Xd_0__inst_mult_5_520 ;
wire Xd_0__inst_mult_5_524 ;
wire Xd_0__inst_mult_5_525 ;
wire Xd_0__inst_mult_5_526 ;
wire Xd_0__inst_mult_5_528 ;
wire Xd_0__inst_mult_5_529 ;
wire Xd_0__inst_mult_5_530 ;
wire Xd_0__inst_mult_5_532 ;
wire Xd_0__inst_mult_5_533 ;
wire Xd_0__inst_mult_5_534 ;
wire Xd_0__inst_mult_2_524 ;
wire Xd_0__inst_mult_2_528 ;
wire Xd_0__inst_mult_2_529 ;
wire Xd_0__inst_mult_2_530 ;
wire Xd_0__inst_mult_2_532 ;
wire Xd_0__inst_mult_2_533 ;
wire Xd_0__inst_mult_2_534 ;
wire Xd_0__inst_mult_2_536 ;
wire Xd_0__inst_mult_2_537 ;
wire Xd_0__inst_mult_2_538 ;
wire Xd_0__inst_mult_3_520 ;
wire Xd_0__inst_mult_3_524 ;
wire Xd_0__inst_mult_3_525 ;
wire Xd_0__inst_mult_3_526 ;
wire Xd_0__inst_mult_3_528 ;
wire Xd_0__inst_mult_3_529 ;
wire Xd_0__inst_mult_3_530 ;
wire Xd_0__inst_mult_3_532 ;
wire Xd_0__inst_mult_3_533 ;
wire Xd_0__inst_mult_3_534 ;
wire Xd_0__inst_mult_0_524 ;
wire Xd_0__inst_mult_0_528 ;
wire Xd_0__inst_mult_0_529 ;
wire Xd_0__inst_mult_0_530 ;
wire Xd_0__inst_mult_0_532 ;
wire Xd_0__inst_mult_0_533 ;
wire Xd_0__inst_mult_0_534 ;
wire Xd_0__inst_mult_0_536 ;
wire Xd_0__inst_mult_0_537 ;
wire Xd_0__inst_mult_0_538 ;
wire Xd_0__inst_mult_1_524 ;
wire Xd_0__inst_mult_1_528 ;
wire Xd_0__inst_mult_1_529 ;
wire Xd_0__inst_mult_1_530 ;
wire Xd_0__inst_mult_1_532 ;
wire Xd_0__inst_mult_1_533 ;
wire Xd_0__inst_mult_1_534 ;
wire Xd_0__inst_mult_1_536 ;
wire Xd_0__inst_mult_1_537 ;
wire Xd_0__inst_mult_1_538 ;
wire Xd_0__inst_mult_12_556 ;
wire Xd_0__inst_mult_12_557 ;
wire Xd_0__inst_mult_12_558 ;
wire Xd_0__inst_mult_14_540 ;
wire Xd_0__inst_mult_14_541 ;
wire Xd_0__inst_mult_14_542 ;
wire Xd_0__inst_mult_13_540 ;
wire Xd_0__inst_mult_13_541 ;
wire Xd_0__inst_mult_13_542 ;
wire Xd_0__inst_mult_13_544 ;
wire Xd_0__inst_mult_13_545 ;
wire Xd_0__inst_mult_13_546 ;
wire Xd_0__inst_mult_1_540 ;
wire Xd_0__inst_mult_1_541 ;
wire Xd_0__inst_mult_1_542 ;
wire Xd_0__inst_mult_14_544 ;
wire Xd_0__inst_mult_14_545 ;
wire Xd_0__inst_mult_14_546 ;
wire Xd_0__inst_mult_14_548 ;
wire Xd_0__inst_mult_14_549 ;
wire Xd_0__inst_mult_14_550 ;
wire Xd_0__inst_mult_15_560 ;
wire Xd_0__inst_mult_15_561 ;
wire Xd_0__inst_mult_15_562 ;
wire Xd_0__inst_mult_15_564 ;
wire Xd_0__inst_mult_15_565 ;
wire Xd_0__inst_mult_15_566 ;
wire Xd_0__inst_mult_14_552 ;
wire Xd_0__inst_mult_14_553 ;
wire Xd_0__inst_mult_14_554 ;
wire Xd_0__inst_mult_10_536 ;
wire Xd_0__inst_mult_10_537 ;
wire Xd_0__inst_mult_10_538 ;
wire Xd_0__inst_mult_10_540 ;
wire Xd_0__inst_mult_10_541 ;
wire Xd_0__inst_mult_10_542 ;
wire Xd_0__inst_mult_0_540 ;
wire Xd_0__inst_mult_0_541 ;
wire Xd_0__inst_mult_0_542 ;
wire Xd_0__inst_mult_11_540 ;
wire Xd_0__inst_mult_11_541 ;
wire Xd_0__inst_mult_11_542 ;
wire Xd_0__inst_mult_11_544 ;
wire Xd_0__inst_mult_11_545 ;
wire Xd_0__inst_mult_11_546 ;
wire Xd_0__inst_mult_3_536 ;
wire Xd_0__inst_mult_3_537 ;
wire Xd_0__inst_mult_3_538 ;
wire Xd_0__inst_mult_8_540 ;
wire Xd_0__inst_mult_8_541 ;
wire Xd_0__inst_mult_8_542 ;
wire Xd_0__inst_mult_8_544 ;
wire Xd_0__inst_mult_8_545 ;
wire Xd_0__inst_mult_8_546 ;
wire Xd_0__inst_mult_2_540 ;
wire Xd_0__inst_mult_2_541 ;
wire Xd_0__inst_mult_2_542 ;
wire Xd_0__inst_mult_9_536 ;
wire Xd_0__inst_mult_9_537 ;
wire Xd_0__inst_mult_9_538 ;
wire Xd_0__inst_mult_9_540 ;
wire Xd_0__inst_mult_9_541 ;
wire Xd_0__inst_mult_9_542 ;
wire Xd_0__inst_mult_1_544 ;
wire Xd_0__inst_mult_1_545 ;
wire Xd_0__inst_mult_1_546 ;
wire Xd_0__inst_mult_6_536 ;
wire Xd_0__inst_mult_6_537 ;
wire Xd_0__inst_mult_6_538 ;
wire Xd_0__inst_mult_6_540 ;
wire Xd_0__inst_mult_6_541 ;
wire Xd_0__inst_mult_6_542 ;
wire Xd_0__inst_mult_5_536 ;
wire Xd_0__inst_mult_5_537 ;
wire Xd_0__inst_mult_5_538 ;
wire Xd_0__inst_mult_7_536 ;
wire Xd_0__inst_mult_7_537 ;
wire Xd_0__inst_mult_7_538 ;
wire Xd_0__inst_mult_7_540 ;
wire Xd_0__inst_mult_7_541 ;
wire Xd_0__inst_mult_7_542 ;
wire Xd_0__inst_mult_7_544 ;
wire Xd_0__inst_mult_7_545 ;
wire Xd_0__inst_mult_7_546 ;
wire Xd_0__inst_mult_4_560 ;
wire Xd_0__inst_mult_4_561 ;
wire Xd_0__inst_mult_4_562 ;
wire Xd_0__inst_mult_6_544 ;
wire Xd_0__inst_mult_6_545 ;
wire Xd_0__inst_mult_6_546 ;
wire Xd_0__inst_mult_5_540 ;
wire Xd_0__inst_mult_5_541 ;
wire Xd_0__inst_mult_5_542 ;
wire Xd_0__inst_mult_5_544 ;
wire Xd_0__inst_mult_5_545 ;
wire Xd_0__inst_mult_5_546 ;
wire Xd_0__inst_mult_9_544 ;
wire Xd_0__inst_mult_9_545 ;
wire Xd_0__inst_mult_9_546 ;
wire Xd_0__inst_mult_2_544 ;
wire Xd_0__inst_mult_2_545 ;
wire Xd_0__inst_mult_2_546 ;
wire Xd_0__inst_mult_2_548 ;
wire Xd_0__inst_mult_2_549 ;
wire Xd_0__inst_mult_2_550 ;
wire Xd_0__inst_mult_13_548 ;
wire Xd_0__inst_mult_13_549 ;
wire Xd_0__inst_mult_13_550 ;
wire Xd_0__inst_mult_3_540 ;
wire Xd_0__inst_mult_3_541 ;
wire Xd_0__inst_mult_3_542 ;
wire Xd_0__inst_mult_3_544 ;
wire Xd_0__inst_mult_3_545 ;
wire Xd_0__inst_mult_3_546 ;
wire Xd_0__inst_mult_8_548 ;
wire Xd_0__inst_mult_8_549 ;
wire Xd_0__inst_mult_8_550 ;
wire Xd_0__inst_mult_0_544 ;
wire Xd_0__inst_mult_0_545 ;
wire Xd_0__inst_mult_0_546 ;
wire Xd_0__inst_mult_0_548 ;
wire Xd_0__inst_mult_0_549 ;
wire Xd_0__inst_mult_0_550 ;
wire Xd_0__inst_mult_11_548 ;
wire Xd_0__inst_mult_11_549 ;
wire Xd_0__inst_mult_11_550 ;
wire Xd_0__inst_mult_1_548 ;
wire Xd_0__inst_mult_1_549 ;
wire Xd_0__inst_mult_1_550 ;
wire Xd_0__inst_mult_1_552 ;
wire Xd_0__inst_mult_1_553 ;
wire Xd_0__inst_mult_1_554 ;
wire Xd_0__inst_mult_10_544 ;
wire Xd_0__inst_mult_10_545 ;
wire Xd_0__inst_mult_10_546 ;
wire Xd_0__inst_mult_12_560 ;
wire Xd_0__inst_mult_12_561 ;
wire Xd_0__inst_mult_12_562 ;
wire Xd_0__inst_mult_13_552 ;
wire Xd_0__inst_mult_13_553 ;
wire Xd_0__inst_mult_13_554 ;
wire Xd_0__inst_mult_13_556 ;
wire Xd_0__inst_mult_13_557 ;
wire Xd_0__inst_mult_13_558 ;
wire Xd_0__inst_mult_14_556 ;
wire Xd_0__inst_mult_14_557 ;
wire Xd_0__inst_mult_14_558 ;
wire Xd_0__inst_mult_14_560 ;
wire Xd_0__inst_mult_14_561 ;
wire Xd_0__inst_mult_14_562 ;
wire Xd_0__inst_mult_15_568 ;
wire Xd_0__inst_mult_15_569 ;
wire Xd_0__inst_mult_15_570 ;
wire Xd_0__inst_mult_10_548 ;
wire Xd_0__inst_mult_10_549 ;
wire Xd_0__inst_mult_10_550 ;
wire Xd_0__inst_mult_10_552 ;
wire Xd_0__inst_mult_10_553 ;
wire Xd_0__inst_mult_10_554 ;
wire Xd_0__inst_mult_11_552 ;
wire Xd_0__inst_mult_11_553 ;
wire Xd_0__inst_mult_11_554 ;
wire Xd_0__inst_mult_11_556 ;
wire Xd_0__inst_mult_11_557 ;
wire Xd_0__inst_mult_11_558 ;
wire Xd_0__inst_mult_8_552 ;
wire Xd_0__inst_mult_8_553 ;
wire Xd_0__inst_mult_8_554 ;
wire Xd_0__inst_mult_8_556 ;
wire Xd_0__inst_mult_8_557 ;
wire Xd_0__inst_mult_8_558 ;
wire Xd_0__inst_mult_9_548 ;
wire Xd_0__inst_mult_9_549 ;
wire Xd_0__inst_mult_9_550 ;
wire Xd_0__inst_mult_9_552 ;
wire Xd_0__inst_mult_9_553 ;
wire Xd_0__inst_mult_9_554 ;
wire Xd_0__inst_mult_6_548 ;
wire Xd_0__inst_mult_6_549 ;
wire Xd_0__inst_mult_6_550 ;
wire Xd_0__inst_mult_6_552 ;
wire Xd_0__inst_mult_6_553 ;
wire Xd_0__inst_mult_6_554 ;
wire Xd_0__inst_mult_7_548 ;
wire Xd_0__inst_mult_7_549 ;
wire Xd_0__inst_mult_7_550 ;
wire Xd_0__inst_mult_7_552 ;
wire Xd_0__inst_mult_7_553 ;
wire Xd_0__inst_mult_7_554 ;
wire Xd_0__inst_mult_4_564 ;
wire Xd_0__inst_mult_4_565 ;
wire Xd_0__inst_mult_4_566 ;
wire Xd_0__inst_mult_5_548 ;
wire Xd_0__inst_mult_5_549 ;
wire Xd_0__inst_mult_5_550 ;
wire Xd_0__inst_mult_5_552 ;
wire Xd_0__inst_mult_5_553 ;
wire Xd_0__inst_mult_5_554 ;
wire Xd_0__inst_mult_2_552 ;
wire Xd_0__inst_mult_2_553 ;
wire Xd_0__inst_mult_2_554 ;
wire Xd_0__inst_mult_2_556 ;
wire Xd_0__inst_mult_2_557 ;
wire Xd_0__inst_mult_2_558 ;
wire Xd_0__inst_mult_3_548 ;
wire Xd_0__inst_mult_3_549 ;
wire Xd_0__inst_mult_3_550 ;
wire Xd_0__inst_mult_3_552 ;
wire Xd_0__inst_mult_3_553 ;
wire Xd_0__inst_mult_3_554 ;
wire Xd_0__inst_mult_0_552 ;
wire Xd_0__inst_mult_0_553 ;
wire Xd_0__inst_mult_0_554 ;
wire Xd_0__inst_mult_0_556 ;
wire Xd_0__inst_mult_0_557 ;
wire Xd_0__inst_mult_0_558 ;
wire Xd_0__inst_mult_1_556 ;
wire Xd_0__inst_mult_1_557 ;
wire Xd_0__inst_mult_1_558 ;
wire Xd_0__inst_mult_1_560 ;
wire Xd_0__inst_mult_1_561 ;
wire Xd_0__inst_mult_1_562 ;
wire Xd_0__inst_mult_12_564 ;
wire Xd_0__inst_mult_13_560 ;
wire Xd_0__inst_mult_13_564 ;
wire Xd_0__inst_mult_13_565 ;
wire Xd_0__inst_mult_13_566 ;
wire Xd_0__inst_mult_14_564 ;
wire Xd_0__inst_mult_14_568 ;
wire Xd_0__inst_mult_14_569 ;
wire Xd_0__inst_mult_14_570 ;
wire Xd_0__inst_mult_15_572 ;
wire Xd_0__inst_mult_10_556 ;
wire Xd_0__inst_mult_10_560 ;
wire Xd_0__inst_mult_10_561 ;
wire Xd_0__inst_mult_10_562 ;
wire Xd_0__inst_mult_11_560 ;
wire Xd_0__inst_mult_11_564 ;
wire Xd_0__inst_mult_11_565 ;
wire Xd_0__inst_mult_11_566 ;
wire Xd_0__inst_mult_8_560 ;
wire Xd_0__inst_mult_8_564 ;
wire Xd_0__inst_mult_8_565 ;
wire Xd_0__inst_mult_8_566 ;
wire Xd_0__inst_mult_9_556 ;
wire Xd_0__inst_mult_9_560 ;
wire Xd_0__inst_mult_9_561 ;
wire Xd_0__inst_mult_9_562 ;
wire Xd_0__inst_mult_6_556 ;
wire Xd_0__inst_mult_6_560 ;
wire Xd_0__inst_mult_6_561 ;
wire Xd_0__inst_mult_6_562 ;
wire Xd_0__inst_mult_7_556 ;
wire Xd_0__inst_mult_7_560 ;
wire Xd_0__inst_mult_7_561 ;
wire Xd_0__inst_mult_7_562 ;
wire Xd_0__inst_mult_4_568 ;
wire Xd_0__inst_mult_5_556 ;
wire Xd_0__inst_mult_5_560 ;
wire Xd_0__inst_mult_5_561 ;
wire Xd_0__inst_mult_5_562 ;
wire Xd_0__inst_mult_2_560 ;
wire Xd_0__inst_mult_2_564 ;
wire Xd_0__inst_mult_2_565 ;
wire Xd_0__inst_mult_2_566 ;
wire Xd_0__inst_mult_3_556 ;
wire Xd_0__inst_mult_3_560 ;
wire Xd_0__inst_mult_3_561 ;
wire Xd_0__inst_mult_3_562 ;
wire Xd_0__inst_mult_0_560 ;
wire Xd_0__inst_mult_0_564 ;
wire Xd_0__inst_mult_0_565 ;
wire Xd_0__inst_mult_0_566 ;
wire Xd_0__inst_mult_1_564 ;
wire Xd_0__inst_mult_1_568 ;
wire Xd_0__inst_mult_1_569 ;
wire Xd_0__inst_mult_1_570 ;
wire Xd_0__inst_mult_13_568 ;
wire Xd_0__inst_mult_13_569 ;
wire Xd_0__inst_mult_13_570 ;
wire Xd_0__inst_mult_14_572 ;
wire Xd_0__inst_mult_14_573 ;
wire Xd_0__inst_mult_14_574 ;
wire Xd_0__inst_mult_10_564 ;
wire Xd_0__inst_mult_10_565 ;
wire Xd_0__inst_mult_10_566 ;
wire Xd_0__inst_mult_11_568 ;
wire Xd_0__inst_mult_11_569 ;
wire Xd_0__inst_mult_11_570 ;
wire Xd_0__inst_mult_8_568 ;
wire Xd_0__inst_mult_8_569 ;
wire Xd_0__inst_mult_8_570 ;
wire Xd_0__inst_mult_9_564 ;
wire Xd_0__inst_mult_9_565 ;
wire Xd_0__inst_mult_9_566 ;
wire Xd_0__inst_mult_6_564 ;
wire Xd_0__inst_mult_6_565 ;
wire Xd_0__inst_mult_6_566 ;
wire Xd_0__inst_mult_7_564 ;
wire Xd_0__inst_mult_7_565 ;
wire Xd_0__inst_mult_7_566 ;
wire Xd_0__inst_mult_5_564 ;
wire Xd_0__inst_mult_5_565 ;
wire Xd_0__inst_mult_5_566 ;
wire Xd_0__inst_mult_2_568 ;
wire Xd_0__inst_mult_2_569 ;
wire Xd_0__inst_mult_2_570 ;
wire Xd_0__inst_mult_3_564 ;
wire Xd_0__inst_mult_3_565 ;
wire Xd_0__inst_mult_3_566 ;
wire Xd_0__inst_mult_0_568 ;
wire Xd_0__inst_mult_0_569 ;
wire Xd_0__inst_mult_0_570 ;
wire Xd_0__inst_mult_1_572 ;
wire Xd_0__inst_mult_1_573 ;
wire Xd_0__inst_mult_1_574 ;
wire Xd_0__inst_mult_13_572 ;
wire Xd_0__inst_mult_14_576 ;
wire Xd_0__inst_mult_10_568 ;
wire Xd_0__inst_mult_11_572 ;
wire Xd_0__inst_mult_8_572 ;
wire Xd_0__inst_mult_9_568 ;
wire Xd_0__inst_mult_6_568 ;
wire Xd_0__inst_mult_7_568 ;
wire Xd_0__inst_mult_5_568 ;
wire Xd_0__inst_mult_2_572 ;
wire Xd_0__inst_mult_3_568 ;
wire Xd_0__inst_mult_0_572 ;
wire Xd_0__inst_mult_1_576 ;
wire Xd_0__inst_mult_12_569 ;
wire Xd_0__inst_mult_12_570 ;
wire Xd_0__inst_mult_13_577 ;
wire Xd_0__inst_mult_13_578 ;
wire Xd_0__inst_mult_10_573 ;
wire Xd_0__inst_mult_10_574 ;
wire Xd_0__inst_mult_11_577 ;
wire Xd_0__inst_mult_11_578 ;
wire Xd_0__inst_mult_8_577 ;
wire Xd_0__inst_mult_8_578 ;
wire Xd_0__inst_mult_9_573 ;
wire Xd_0__inst_mult_9_574 ;
wire Xd_0__inst_mult_6_573 ;
wire Xd_0__inst_mult_6_574 ;
wire Xd_0__inst_mult_7_573 ;
wire Xd_0__inst_mult_7_574 ;
wire Xd_0__inst_mult_4_573 ;
wire Xd_0__inst_mult_4_574 ;
wire Xd_0__inst_mult_5_573 ;
wire Xd_0__inst_mult_5_574 ;
wire Xd_0__inst_mult_2_577 ;
wire Xd_0__inst_mult_2_578 ;
wire Xd_0__inst_mult_3_573 ;
wire Xd_0__inst_mult_3_574 ;
wire Xd_0__inst_mult_0_577 ;
wire Xd_0__inst_mult_0_578 ;
wire Xd_0__inst_mult_12_573 ;
wire Xd_0__inst_mult_12_574 ;
wire Xd_0__inst_mult_13_581 ;
wire Xd_0__inst_mult_13_582 ;
wire Xd_0__inst_mult_14_581 ;
wire Xd_0__inst_mult_14_582 ;
wire Xd_0__inst_mult_15_577 ;
wire Xd_0__inst_mult_15_578 ;
wire Xd_0__inst_mult_10_577 ;
wire Xd_0__inst_mult_10_578 ;
wire Xd_0__inst_mult_11_581 ;
wire Xd_0__inst_mult_11_582 ;
wire Xd_0__inst_mult_8_581 ;
wire Xd_0__inst_mult_8_582 ;
wire Xd_0__inst_mult_9_577 ;
wire Xd_0__inst_mult_9_578 ;
wire Xd_0__inst_mult_6_577 ;
wire Xd_0__inst_mult_6_578 ;
wire Xd_0__inst_mult_7_577 ;
wire Xd_0__inst_mult_7_578 ;
wire Xd_0__inst_mult_4_577 ;
wire Xd_0__inst_mult_4_578 ;
wire Xd_0__inst_mult_5_577 ;
wire Xd_0__inst_mult_5_578 ;
wire Xd_0__inst_mult_2_581 ;
wire Xd_0__inst_mult_2_582 ;
wire Xd_0__inst_mult_3_577 ;
wire Xd_0__inst_mult_3_578 ;
wire Xd_0__inst_mult_0_581 ;
wire Xd_0__inst_mult_0_582 ;
wire Xd_0__inst_mult_1_581 ;
wire Xd_0__inst_mult_1_582 ;
wire Xd_0__inst_mult_12_577 ;
wire Xd_0__inst_mult_12_578 ;
wire Xd_0__inst_mult_13_585 ;
wire Xd_0__inst_mult_13_586 ;
wire Xd_0__inst_mult_14_585 ;
wire Xd_0__inst_mult_14_586 ;
wire Xd_0__inst_mult_15_581 ;
wire Xd_0__inst_mult_15_582 ;
wire Xd_0__inst_mult_10_581 ;
wire Xd_0__inst_mult_10_582 ;
wire Xd_0__inst_mult_11_585 ;
wire Xd_0__inst_mult_11_586 ;
wire Xd_0__inst_mult_8_585 ;
wire Xd_0__inst_mult_8_586 ;
wire Xd_0__inst_mult_9_581 ;
wire Xd_0__inst_mult_9_582 ;
wire Xd_0__inst_mult_6_581 ;
wire Xd_0__inst_mult_6_582 ;
wire Xd_0__inst_mult_7_581 ;
wire Xd_0__inst_mult_7_582 ;
wire Xd_0__inst_mult_4_581 ;
wire Xd_0__inst_mult_4_582 ;
wire Xd_0__inst_mult_5_581 ;
wire Xd_0__inst_mult_5_582 ;
wire Xd_0__inst_mult_2_585 ;
wire Xd_0__inst_mult_2_586 ;
wire Xd_0__inst_mult_3_581 ;
wire Xd_0__inst_mult_3_582 ;
wire Xd_0__inst_mult_0_585 ;
wire Xd_0__inst_mult_0_586 ;
wire Xd_0__inst_mult_1_585 ;
wire Xd_0__inst_mult_1_586 ;
wire Xd_0__inst_mult_12_581 ;
wire Xd_0__inst_mult_12_582 ;
wire Xd_0__inst_mult_15_585 ;
wire Xd_0__inst_mult_15_586 ;
wire Xd_0__inst_mult_4_585 ;
wire Xd_0__inst_mult_4_586 ;
wire Xd_0__inst_inst_first_level_2__0__q ;
wire Xd_0__inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_first_level_2__1__q ;
wire Xd_0__inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_first_level_2__2__q ;
wire Xd_0__inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_first_level_2__3__q ;
wire Xd_0__inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_first_level_2__4__q ;
wire Xd_0__inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_first_level_2__5__q ;
wire Xd_0__inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_first_level_2__6__q ;
wire Xd_0__inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_first_level_2__7__q ;
wire Xd_0__inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_first_level_2__8__q ;
wire Xd_0__inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_first_level_2__9__q ;
wire Xd_0__inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_first_level_2__10__q ;
wire Xd_0__inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_first_level_2__11__q ;
wire Xd_0__inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_first_level_2__12__q ;
wire Xd_0__inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_first_level_2__13__q ;
wire Xd_0__inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_first_level_2__14__q ;
wire Xd_0__inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_first_level_2__15__q ;
wire Xd_0__inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_first_level_2__16__q ;
wire Xd_0__inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_first_level_2__17__q ;
wire Xd_0__inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_first_level_0__17__q ;
wire Xd_0__inst_inst_first_level_2__18__q ;
wire Xd_0__inst_inst_first_level_1__18__q ;
wire Xd_0__inst_inst_first_level_0__18__q ;
wire Xd_0__inst_inst_first_level_2__19__q ;
wire Xd_0__inst_inst_first_level_1__19__q ;
wire Xd_0__inst_inst_first_level_0__19__q ;
wire Xd_0__inst_inst_first_level_2__20__q ;
wire Xd_0__inst_inst_first_level_1__20__q ;
wire Xd_0__inst_inst_first_level_0__20__q ;
wire Xd_0__inst_inst_first_level_2__21__q ;
wire Xd_0__inst_inst_first_level_1__21__q ;
wire Xd_0__inst_inst_first_level_0__21__q ;
wire Xd_0__inst_inst_first_level_2__22__q ;
wire Xd_0__inst_inst_first_level_1__22__q ;
wire Xd_0__inst_inst_first_level_0__22__q ;
wire Xd_0__inst_inst_first_level_2__23__q ;
wire Xd_0__inst_inst_first_level_1__23__q ;
wire Xd_0__inst_inst_first_level_0__23__q ;
wire Xd_0__inst_inst_first_level_2__25__q ;
wire Xd_0__inst_inst_first_level_1__24__q ;
wire Xd_0__inst_inst_first_level_0__24__q ;
wire Xd_0__inst_inst_first_level_1__25__q ;
wire Xd_0__inst_inst_first_level_0__25__q ;
wire Xd_0__inst_r_sum1_6__0__q ;
wire Xd_0__inst_r_sum1_7__0__q ;
wire Xd_0__inst_r_sum1_5__0__q ;
wire Xd_0__inst_r_sum1_4__0__q ;
wire Xd_0__inst_r_sum1_3__0__q ;
wire Xd_0__inst_r_sum1_2__0__q ;
wire Xd_0__inst_r_sum1_1__0__q ;
wire Xd_0__inst_r_sum1_0__0__q ;
wire Xd_0__inst_r_sum1_6__1__q ;
wire Xd_0__inst_r_sum1_7__1__q ;
wire Xd_0__inst_r_sum1_5__1__q ;
wire Xd_0__inst_r_sum1_4__1__q ;
wire Xd_0__inst_r_sum1_3__1__q ;
wire Xd_0__inst_r_sum1_2__1__q ;
wire Xd_0__inst_r_sum1_1__1__q ;
wire Xd_0__inst_r_sum1_0__1__q ;
wire Xd_0__inst_r_sum1_6__2__q ;
wire Xd_0__inst_r_sum1_7__2__q ;
wire Xd_0__inst_r_sum1_5__2__q ;
wire Xd_0__inst_r_sum1_4__2__q ;
wire Xd_0__inst_r_sum1_3__2__q ;
wire Xd_0__inst_r_sum1_2__2__q ;
wire Xd_0__inst_r_sum1_1__2__q ;
wire Xd_0__inst_r_sum1_0__2__q ;
wire Xd_0__inst_r_sum1_6__3__q ;
wire Xd_0__inst_r_sum1_7__3__q ;
wire Xd_0__inst_r_sum1_5__3__q ;
wire Xd_0__inst_r_sum1_4__3__q ;
wire Xd_0__inst_r_sum1_3__3__q ;
wire Xd_0__inst_r_sum1_2__3__q ;
wire Xd_0__inst_r_sum1_1__3__q ;
wire Xd_0__inst_r_sum1_0__3__q ;
wire Xd_0__inst_r_sum1_6__4__q ;
wire Xd_0__inst_r_sum1_7__4__q ;
wire Xd_0__inst_r_sum1_5__4__q ;
wire Xd_0__inst_r_sum1_4__4__q ;
wire Xd_0__inst_r_sum1_3__4__q ;
wire Xd_0__inst_r_sum1_2__4__q ;
wire Xd_0__inst_r_sum1_1__4__q ;
wire Xd_0__inst_r_sum1_0__4__q ;
wire Xd_0__inst_r_sum1_6__5__q ;
wire Xd_0__inst_r_sum1_7__5__q ;
wire Xd_0__inst_r_sum1_5__5__q ;
wire Xd_0__inst_r_sum1_4__5__q ;
wire Xd_0__inst_r_sum1_3__5__q ;
wire Xd_0__inst_r_sum1_2__5__q ;
wire Xd_0__inst_r_sum1_1__5__q ;
wire Xd_0__inst_r_sum1_0__5__q ;
wire Xd_0__inst_r_sum1_6__6__q ;
wire Xd_0__inst_r_sum1_7__6__q ;
wire Xd_0__inst_r_sum1_5__6__q ;
wire Xd_0__inst_r_sum1_4__6__q ;
wire Xd_0__inst_r_sum1_3__6__q ;
wire Xd_0__inst_r_sum1_2__6__q ;
wire Xd_0__inst_r_sum1_1__6__q ;
wire Xd_0__inst_r_sum1_0__6__q ;
wire Xd_0__inst_r_sum1_6__7__q ;
wire Xd_0__inst_r_sum1_7__7__q ;
wire Xd_0__inst_r_sum1_5__7__q ;
wire Xd_0__inst_r_sum1_4__7__q ;
wire Xd_0__inst_r_sum1_3__7__q ;
wire Xd_0__inst_r_sum1_2__7__q ;
wire Xd_0__inst_r_sum1_1__7__q ;
wire Xd_0__inst_r_sum1_0__7__q ;
wire Xd_0__inst_r_sum1_6__8__q ;
wire Xd_0__inst_r_sum1_7__8__q ;
wire Xd_0__inst_r_sum1_5__8__q ;
wire Xd_0__inst_r_sum1_4__8__q ;
wire Xd_0__inst_r_sum1_3__8__q ;
wire Xd_0__inst_r_sum1_2__8__q ;
wire Xd_0__inst_r_sum1_1__8__q ;
wire Xd_0__inst_r_sum1_0__8__q ;
wire Xd_0__inst_r_sum1_6__9__q ;
wire Xd_0__inst_r_sum1_7__9__q ;
wire Xd_0__inst_r_sum1_5__9__q ;
wire Xd_0__inst_r_sum1_4__9__q ;
wire Xd_0__inst_r_sum1_3__9__q ;
wire Xd_0__inst_r_sum1_2__9__q ;
wire Xd_0__inst_r_sum1_1__9__q ;
wire Xd_0__inst_r_sum1_0__9__q ;
wire Xd_0__inst_r_sum1_6__10__q ;
wire Xd_0__inst_r_sum1_7__10__q ;
wire Xd_0__inst_r_sum1_5__10__q ;
wire Xd_0__inst_r_sum1_4__10__q ;
wire Xd_0__inst_r_sum1_3__10__q ;
wire Xd_0__inst_r_sum1_2__10__q ;
wire Xd_0__inst_r_sum1_1__10__q ;
wire Xd_0__inst_r_sum1_0__10__q ;
wire Xd_0__inst_r_sum1_6__11__q ;
wire Xd_0__inst_r_sum1_7__11__q ;
wire Xd_0__inst_r_sum1_5__11__q ;
wire Xd_0__inst_r_sum1_4__11__q ;
wire Xd_0__inst_r_sum1_3__11__q ;
wire Xd_0__inst_r_sum1_2__11__q ;
wire Xd_0__inst_r_sum1_1__11__q ;
wire Xd_0__inst_r_sum1_0__11__q ;
wire Xd_0__inst_r_sum1_6__12__q ;
wire Xd_0__inst_r_sum1_7__12__q ;
wire Xd_0__inst_r_sum1_5__12__q ;
wire Xd_0__inst_r_sum1_4__12__q ;
wire Xd_0__inst_r_sum1_3__12__q ;
wire Xd_0__inst_r_sum1_2__12__q ;
wire Xd_0__inst_r_sum1_1__12__q ;
wire Xd_0__inst_r_sum1_0__12__q ;
wire Xd_0__inst_r_sum1_6__13__q ;
wire Xd_0__inst_r_sum1_7__13__q ;
wire Xd_0__inst_r_sum1_5__13__q ;
wire Xd_0__inst_r_sum1_4__13__q ;
wire Xd_0__inst_r_sum1_3__13__q ;
wire Xd_0__inst_r_sum1_2__13__q ;
wire Xd_0__inst_r_sum1_1__13__q ;
wire Xd_0__inst_r_sum1_0__13__q ;
wire Xd_0__inst_r_sum1_6__14__q ;
wire Xd_0__inst_r_sum1_7__14__q ;
wire Xd_0__inst_r_sum1_5__14__q ;
wire Xd_0__inst_r_sum1_4__14__q ;
wire Xd_0__inst_r_sum1_3__14__q ;
wire Xd_0__inst_r_sum1_2__14__q ;
wire Xd_0__inst_r_sum1_1__14__q ;
wire Xd_0__inst_r_sum1_0__14__q ;
wire Xd_0__inst_r_sum1_6__15__q ;
wire Xd_0__inst_r_sum1_7__15__q ;
wire Xd_0__inst_r_sum1_5__15__q ;
wire Xd_0__inst_r_sum1_4__15__q ;
wire Xd_0__inst_r_sum1_3__15__q ;
wire Xd_0__inst_r_sum1_2__15__q ;
wire Xd_0__inst_r_sum1_1__15__q ;
wire Xd_0__inst_r_sum1_0__15__q ;
wire Xd_0__inst_r_sum1_6__16__q ;
wire Xd_0__inst_r_sum1_7__16__q ;
wire Xd_0__inst_r_sum1_5__16__q ;
wire Xd_0__inst_r_sum1_4__16__q ;
wire Xd_0__inst_r_sum1_3__16__q ;
wire Xd_0__inst_r_sum1_2__16__q ;
wire Xd_0__inst_r_sum1_1__16__q ;
wire Xd_0__inst_r_sum1_0__16__q ;
wire Xd_0__inst_r_sum1_6__17__q ;
wire Xd_0__inst_r_sum1_7__17__q ;
wire Xd_0__inst_r_sum1_5__17__q ;
wire Xd_0__inst_r_sum1_4__17__q ;
wire Xd_0__inst_r_sum1_3__17__q ;
wire Xd_0__inst_r_sum1_2__17__q ;
wire Xd_0__inst_r_sum1_1__17__q ;
wire Xd_0__inst_r_sum1_0__17__q ;
wire Xd_0__inst_r_sum1_6__18__q ;
wire Xd_0__inst_r_sum1_7__18__q ;
wire Xd_0__inst_r_sum1_5__18__q ;
wire Xd_0__inst_r_sum1_4__18__q ;
wire Xd_0__inst_r_sum1_3__18__q ;
wire Xd_0__inst_r_sum1_2__18__q ;
wire Xd_0__inst_r_sum1_1__18__q ;
wire Xd_0__inst_r_sum1_0__18__q ;
wire Xd_0__inst_r_sum1_6__19__q ;
wire Xd_0__inst_r_sum1_7__19__q ;
wire Xd_0__inst_r_sum1_5__19__q ;
wire Xd_0__inst_r_sum1_4__19__q ;
wire Xd_0__inst_r_sum1_3__19__q ;
wire Xd_0__inst_r_sum1_2__19__q ;
wire Xd_0__inst_r_sum1_1__19__q ;
wire Xd_0__inst_r_sum1_0__19__q ;
wire Xd_0__inst_r_sum1_6__20__q ;
wire Xd_0__inst_r_sum1_7__20__q ;
wire Xd_0__inst_r_sum1_5__20__q ;
wire Xd_0__inst_r_sum1_4__20__q ;
wire Xd_0__inst_r_sum1_3__20__q ;
wire Xd_0__inst_r_sum1_2__20__q ;
wire Xd_0__inst_r_sum1_1__20__q ;
wire Xd_0__inst_r_sum1_0__20__q ;
wire Xd_0__inst_r_sum1_6__21__q ;
wire Xd_0__inst_r_sum1_7__21__q ;
wire Xd_0__inst_r_sum1_5__21__q ;
wire Xd_0__inst_r_sum1_4__21__q ;
wire Xd_0__inst_r_sum1_3__21__q ;
wire Xd_0__inst_r_sum1_2__21__q ;
wire Xd_0__inst_r_sum1_1__21__q ;
wire Xd_0__inst_r_sum1_0__21__q ;
wire Xd_0__inst_r_sum1_6__22__q ;
wire Xd_0__inst_r_sum1_7__22__q ;
wire Xd_0__inst_r_sum1_5__22__q ;
wire Xd_0__inst_r_sum1_4__22__q ;
wire Xd_0__inst_r_sum1_3__22__q ;
wire Xd_0__inst_r_sum1_2__22__q ;
wire Xd_0__inst_r_sum1_1__22__q ;
wire Xd_0__inst_r_sum1_0__22__q ;
wire Xd_0__inst_r_sum1_6__23__q ;
wire Xd_0__inst_r_sum1_7__23__q ;
wire Xd_0__inst_r_sum1_5__23__q ;
wire Xd_0__inst_r_sum1_4__23__q ;
wire Xd_0__inst_r_sum1_3__23__q ;
wire Xd_0__inst_r_sum1_2__23__q ;
wire Xd_0__inst_r_sum1_1__23__q ;
wire Xd_0__inst_r_sum1_0__23__q ;
wire Xd_0__inst_product_12__0__q ;
wire Xd_0__inst_product_13__0__q ;
wire Xd_0__inst_product_14__0__q ;
wire Xd_0__inst_product_15__0__q ;
wire Xd_0__inst_product_10__0__q ;
wire Xd_0__inst_product_11__0__q ;
wire Xd_0__inst_product_8__0__q ;
wire Xd_0__inst_product_9__0__q ;
wire Xd_0__inst_product_6__0__q ;
wire Xd_0__inst_product_7__0__q ;
wire Xd_0__inst_product_4__0__q ;
wire Xd_0__inst_product_5__0__q ;
wire Xd_0__inst_product_2__0__q ;
wire Xd_0__inst_product_3__0__q ;
wire Xd_0__inst_product_0__0__q ;
wire Xd_0__inst_product_1__0__q ;
wire Xd_0__inst_product_12__1__q ;
wire Xd_0__inst_product_13__1__q ;
wire Xd_0__inst_product_14__1__q ;
wire Xd_0__inst_product_15__1__q ;
wire Xd_0__inst_product_10__1__q ;
wire Xd_0__inst_product_11__1__q ;
wire Xd_0__inst_product_8__1__q ;
wire Xd_0__inst_product_9__1__q ;
wire Xd_0__inst_product_6__1__q ;
wire Xd_0__inst_product_7__1__q ;
wire Xd_0__inst_product_4__1__q ;
wire Xd_0__inst_product_5__1__q ;
wire Xd_0__inst_product_2__1__q ;
wire Xd_0__inst_product_3__1__q ;
wire Xd_0__inst_product_0__1__q ;
wire Xd_0__inst_product_1__1__q ;
wire Xd_0__inst_product_12__2__q ;
wire Xd_0__inst_product_13__2__q ;
wire Xd_0__inst_product_14__2__q ;
wire Xd_0__inst_product_15__2__q ;
wire Xd_0__inst_product_10__2__q ;
wire Xd_0__inst_product_11__2__q ;
wire Xd_0__inst_product_8__2__q ;
wire Xd_0__inst_product_9__2__q ;
wire Xd_0__inst_product_6__2__q ;
wire Xd_0__inst_product_7__2__q ;
wire Xd_0__inst_product_4__2__q ;
wire Xd_0__inst_product_5__2__q ;
wire Xd_0__inst_product_2__2__q ;
wire Xd_0__inst_product_3__2__q ;
wire Xd_0__inst_product_0__2__q ;
wire Xd_0__inst_product_1__2__q ;
wire Xd_0__inst_product_12__3__q ;
wire Xd_0__inst_product_13__3__q ;
wire Xd_0__inst_product_14__3__q ;
wire Xd_0__inst_product_15__3__q ;
wire Xd_0__inst_product_10__3__q ;
wire Xd_0__inst_product_11__3__q ;
wire Xd_0__inst_product_8__3__q ;
wire Xd_0__inst_product_9__3__q ;
wire Xd_0__inst_product_6__3__q ;
wire Xd_0__inst_product_7__3__q ;
wire Xd_0__inst_product_4__3__q ;
wire Xd_0__inst_product_5__3__q ;
wire Xd_0__inst_product_2__3__q ;
wire Xd_0__inst_product_3__3__q ;
wire Xd_0__inst_product_0__3__q ;
wire Xd_0__inst_product_1__3__q ;
wire Xd_0__inst_product_12__4__q ;
wire Xd_0__inst_product_13__4__q ;
wire Xd_0__inst_product_14__4__q ;
wire Xd_0__inst_product_15__4__q ;
wire Xd_0__inst_product_10__4__q ;
wire Xd_0__inst_product_11__4__q ;
wire Xd_0__inst_product_8__4__q ;
wire Xd_0__inst_product_9__4__q ;
wire Xd_0__inst_product_6__4__q ;
wire Xd_0__inst_product_7__4__q ;
wire Xd_0__inst_product_4__4__q ;
wire Xd_0__inst_product_5__4__q ;
wire Xd_0__inst_product_2__4__q ;
wire Xd_0__inst_product_3__4__q ;
wire Xd_0__inst_product_0__4__q ;
wire Xd_0__inst_product_1__4__q ;
wire Xd_0__inst_product_12__5__q ;
wire Xd_0__inst_product_13__5__q ;
wire Xd_0__inst_product_14__5__q ;
wire Xd_0__inst_product_15__5__q ;
wire Xd_0__inst_product_10__5__q ;
wire Xd_0__inst_product_11__5__q ;
wire Xd_0__inst_product_8__5__q ;
wire Xd_0__inst_product_9__5__q ;
wire Xd_0__inst_product_6__5__q ;
wire Xd_0__inst_product_7__5__q ;
wire Xd_0__inst_product_4__5__q ;
wire Xd_0__inst_product_5__5__q ;
wire Xd_0__inst_product_2__5__q ;
wire Xd_0__inst_product_3__5__q ;
wire Xd_0__inst_product_0__5__q ;
wire Xd_0__inst_product_1__5__q ;
wire Xd_0__inst_product_12__6__q ;
wire Xd_0__inst_product_13__6__q ;
wire Xd_0__inst_product_14__6__q ;
wire Xd_0__inst_product_15__6__q ;
wire Xd_0__inst_product_10__6__q ;
wire Xd_0__inst_product_11__6__q ;
wire Xd_0__inst_product_8__6__q ;
wire Xd_0__inst_product_9__6__q ;
wire Xd_0__inst_product_6__6__q ;
wire Xd_0__inst_product_7__6__q ;
wire Xd_0__inst_product_4__6__q ;
wire Xd_0__inst_product_5__6__q ;
wire Xd_0__inst_product_2__6__q ;
wire Xd_0__inst_product_3__6__q ;
wire Xd_0__inst_product_0__6__q ;
wire Xd_0__inst_product_1__6__q ;
wire Xd_0__inst_product_12__7__q ;
wire Xd_0__inst_product_13__7__q ;
wire Xd_0__inst_product_14__7__q ;
wire Xd_0__inst_product_15__7__q ;
wire Xd_0__inst_product_10__7__q ;
wire Xd_0__inst_product_11__7__q ;
wire Xd_0__inst_product_8__7__q ;
wire Xd_0__inst_product_9__7__q ;
wire Xd_0__inst_product_6__7__q ;
wire Xd_0__inst_product_7__7__q ;
wire Xd_0__inst_product_4__7__q ;
wire Xd_0__inst_product_5__7__q ;
wire Xd_0__inst_product_2__7__q ;
wire Xd_0__inst_product_3__7__q ;
wire Xd_0__inst_product_0__7__q ;
wire Xd_0__inst_product_1__7__q ;
wire Xd_0__inst_product_12__8__q ;
wire Xd_0__inst_product_13__8__q ;
wire Xd_0__inst_product_14__8__q ;
wire Xd_0__inst_product_15__8__q ;
wire Xd_0__inst_product_10__8__q ;
wire Xd_0__inst_product_11__8__q ;
wire Xd_0__inst_product_8__8__q ;
wire Xd_0__inst_product_9__8__q ;
wire Xd_0__inst_product_6__8__q ;
wire Xd_0__inst_product_7__8__q ;
wire Xd_0__inst_product_4__8__q ;
wire Xd_0__inst_product_5__8__q ;
wire Xd_0__inst_product_2__8__q ;
wire Xd_0__inst_product_3__8__q ;
wire Xd_0__inst_product_0__8__q ;
wire Xd_0__inst_product_1__8__q ;
wire Xd_0__inst_product_12__9__q ;
wire Xd_0__inst_product_13__9__q ;
wire Xd_0__inst_product_14__9__q ;
wire Xd_0__inst_product_15__9__q ;
wire Xd_0__inst_product_10__9__q ;
wire Xd_0__inst_product_11__9__q ;
wire Xd_0__inst_product_8__9__q ;
wire Xd_0__inst_product_9__9__q ;
wire Xd_0__inst_product_6__9__q ;
wire Xd_0__inst_product_7__9__q ;
wire Xd_0__inst_product_4__9__q ;
wire Xd_0__inst_product_5__9__q ;
wire Xd_0__inst_product_2__9__q ;
wire Xd_0__inst_product_3__9__q ;
wire Xd_0__inst_product_0__9__q ;
wire Xd_0__inst_product_1__9__q ;
wire Xd_0__inst_product_12__10__q ;
wire Xd_0__inst_product_13__10__q ;
wire Xd_0__inst_product_14__10__q ;
wire Xd_0__inst_product_15__10__q ;
wire Xd_0__inst_product_10__10__q ;
wire Xd_0__inst_product_11__10__q ;
wire Xd_0__inst_product_8__10__q ;
wire Xd_0__inst_product_9__10__q ;
wire Xd_0__inst_product_6__10__q ;
wire Xd_0__inst_product_7__10__q ;
wire Xd_0__inst_product_4__10__q ;
wire Xd_0__inst_product_5__10__q ;
wire Xd_0__inst_product_2__10__q ;
wire Xd_0__inst_product_3__10__q ;
wire Xd_0__inst_product_0__10__q ;
wire Xd_0__inst_product_1__10__q ;
wire Xd_0__inst_product_12__11__q ;
wire Xd_0__inst_product_13__11__q ;
wire Xd_0__inst_product_14__11__q ;
wire Xd_0__inst_product_15__11__q ;
wire Xd_0__inst_product_10__11__q ;
wire Xd_0__inst_product_11__11__q ;
wire Xd_0__inst_product_8__11__q ;
wire Xd_0__inst_product_9__11__q ;
wire Xd_0__inst_product_6__11__q ;
wire Xd_0__inst_product_7__11__q ;
wire Xd_0__inst_product_4__11__q ;
wire Xd_0__inst_product_5__11__q ;
wire Xd_0__inst_product_2__11__q ;
wire Xd_0__inst_product_3__11__q ;
wire Xd_0__inst_product_0__11__q ;
wire Xd_0__inst_product_1__11__q ;
wire Xd_0__inst_product_12__12__q ;
wire Xd_0__inst_product_13__12__q ;
wire Xd_0__inst_product_14__12__q ;
wire Xd_0__inst_product_15__12__q ;
wire Xd_0__inst_product_10__12__q ;
wire Xd_0__inst_product_11__12__q ;
wire Xd_0__inst_product_8__12__q ;
wire Xd_0__inst_product_9__12__q ;
wire Xd_0__inst_product_6__12__q ;
wire Xd_0__inst_product_7__12__q ;
wire Xd_0__inst_product_4__12__q ;
wire Xd_0__inst_product_5__12__q ;
wire Xd_0__inst_product_2__12__q ;
wire Xd_0__inst_product_3__12__q ;
wire Xd_0__inst_product_0__12__q ;
wire Xd_0__inst_product_1__12__q ;
wire Xd_0__inst_product_12__13__q ;
wire Xd_0__inst_product_13__13__q ;
wire Xd_0__inst_product_14__13__q ;
wire Xd_0__inst_product_15__13__q ;
wire Xd_0__inst_product_10__13__q ;
wire Xd_0__inst_product_11__13__q ;
wire Xd_0__inst_product_8__13__q ;
wire Xd_0__inst_product_9__13__q ;
wire Xd_0__inst_product_6__13__q ;
wire Xd_0__inst_product_7__13__q ;
wire Xd_0__inst_product_4__13__q ;
wire Xd_0__inst_product_5__13__q ;
wire Xd_0__inst_product_2__13__q ;
wire Xd_0__inst_product_3__13__q ;
wire Xd_0__inst_product_0__13__q ;
wire Xd_0__inst_product_1__13__q ;
wire Xd_0__inst_product_12__14__q ;
wire Xd_0__inst_product_13__14__q ;
wire Xd_0__inst_product_14__14__q ;
wire Xd_0__inst_product_15__14__q ;
wire Xd_0__inst_product_10__14__q ;
wire Xd_0__inst_product_11__14__q ;
wire Xd_0__inst_product_8__14__q ;
wire Xd_0__inst_product_9__14__q ;
wire Xd_0__inst_product_6__14__q ;
wire Xd_0__inst_product_7__14__q ;
wire Xd_0__inst_product_4__14__q ;
wire Xd_0__inst_product_5__14__q ;
wire Xd_0__inst_product_2__14__q ;
wire Xd_0__inst_product_3__14__q ;
wire Xd_0__inst_product_0__14__q ;
wire Xd_0__inst_product_1__14__q ;
wire Xd_0__inst_product_12__15__q ;
wire Xd_0__inst_product_13__15__q ;
wire Xd_0__inst_product_14__15__q ;
wire Xd_0__inst_product_15__15__q ;
wire Xd_0__inst_product_10__15__q ;
wire Xd_0__inst_product_11__15__q ;
wire Xd_0__inst_product_8__15__q ;
wire Xd_0__inst_product_9__15__q ;
wire Xd_0__inst_product_6__15__q ;
wire Xd_0__inst_product_7__15__q ;
wire Xd_0__inst_product_4__15__q ;
wire Xd_0__inst_product_5__15__q ;
wire Xd_0__inst_product_2__15__q ;
wire Xd_0__inst_product_3__15__q ;
wire Xd_0__inst_product_0__15__q ;
wire Xd_0__inst_product_1__15__q ;
wire Xd_0__inst_product_12__16__q ;
wire Xd_0__inst_product_13__16__q ;
wire Xd_0__inst_product_14__16__q ;
wire Xd_0__inst_product_15__16__q ;
wire Xd_0__inst_product_10__16__q ;
wire Xd_0__inst_product_11__16__q ;
wire Xd_0__inst_product_8__16__q ;
wire Xd_0__inst_product_9__16__q ;
wire Xd_0__inst_product_6__16__q ;
wire Xd_0__inst_product_7__16__q ;
wire Xd_0__inst_product_4__16__q ;
wire Xd_0__inst_product_5__16__q ;
wire Xd_0__inst_product_2__16__q ;
wire Xd_0__inst_product_3__16__q ;
wire Xd_0__inst_product_0__16__q ;
wire Xd_0__inst_product_1__16__q ;
wire Xd_0__inst_product_12__17__q ;
wire Xd_0__inst_product_13__17__q ;
wire Xd_0__inst_product_14__17__q ;
wire Xd_0__inst_product_15__17__q ;
wire Xd_0__inst_product_10__17__q ;
wire Xd_0__inst_product_11__17__q ;
wire Xd_0__inst_product_8__17__q ;
wire Xd_0__inst_product_9__17__q ;
wire Xd_0__inst_product_6__17__q ;
wire Xd_0__inst_product_7__17__q ;
wire Xd_0__inst_product_4__17__q ;
wire Xd_0__inst_product_5__17__q ;
wire Xd_0__inst_product_2__17__q ;
wire Xd_0__inst_product_3__17__q ;
wire Xd_0__inst_product_0__17__q ;
wire Xd_0__inst_product_1__17__q ;
wire Xd_0__inst_product_12__18__q ;
wire Xd_0__inst_product_13__18__q ;
wire Xd_0__inst_product_14__18__q ;
wire Xd_0__inst_product_15__18__q ;
wire Xd_0__inst_product_10__18__q ;
wire Xd_0__inst_product_11__18__q ;
wire Xd_0__inst_product_8__18__q ;
wire Xd_0__inst_product_9__18__q ;
wire Xd_0__inst_product_6__18__q ;
wire Xd_0__inst_product_7__18__q ;
wire Xd_0__inst_product_4__18__q ;
wire Xd_0__inst_product_5__18__q ;
wire Xd_0__inst_product_2__18__q ;
wire Xd_0__inst_product_3__18__q ;
wire Xd_0__inst_product_0__18__q ;
wire Xd_0__inst_product_1__18__q ;
wire Xd_0__inst_product_12__19__q ;
wire Xd_0__inst_product_13__19__q ;
wire Xd_0__inst_product_14__19__q ;
wire Xd_0__inst_product_15__19__q ;
wire Xd_0__inst_product_10__19__q ;
wire Xd_0__inst_product_11__19__q ;
wire Xd_0__inst_product_8__19__q ;
wire Xd_0__inst_product_9__19__q ;
wire Xd_0__inst_product_6__19__q ;
wire Xd_0__inst_product_7__19__q ;
wire Xd_0__inst_product_4__19__q ;
wire Xd_0__inst_product_5__19__q ;
wire Xd_0__inst_product_2__19__q ;
wire Xd_0__inst_product_3__19__q ;
wire Xd_0__inst_product_0__19__q ;
wire Xd_0__inst_product_1__19__q ;
wire Xd_0__inst_product_12__20__q ;
wire Xd_0__inst_product_13__20__q ;
wire Xd_0__inst_product_14__20__q ;
wire Xd_0__inst_product_15__20__q ;
wire Xd_0__inst_product_10__20__q ;
wire Xd_0__inst_product_11__20__q ;
wire Xd_0__inst_product_8__20__q ;
wire Xd_0__inst_product_9__20__q ;
wire Xd_0__inst_product_6__20__q ;
wire Xd_0__inst_product_7__20__q ;
wire Xd_0__inst_product_4__20__q ;
wire Xd_0__inst_product_5__20__q ;
wire Xd_0__inst_product_2__20__q ;
wire Xd_0__inst_product_3__20__q ;
wire Xd_0__inst_product_0__20__q ;
wire Xd_0__inst_product_1__20__q ;
wire Xd_0__inst_product_12__21__q ;
wire Xd_0__inst_product_13__21__q ;
wire Xd_0__inst_product_14__21__q ;
wire Xd_0__inst_product_15__21__q ;
wire Xd_0__inst_product_10__21__q ;
wire Xd_0__inst_product_11__21__q ;
wire Xd_0__inst_product_8__21__q ;
wire Xd_0__inst_product_9__21__q ;
wire Xd_0__inst_product_6__21__q ;
wire Xd_0__inst_product_7__21__q ;
wire Xd_0__inst_product_4__21__q ;
wire Xd_0__inst_product_5__21__q ;
wire Xd_0__inst_product_2__21__q ;
wire Xd_0__inst_product_3__21__q ;
wire Xd_0__inst_product_0__21__q ;
wire Xd_0__inst_product_1__21__q ;
wire Xd_0__inst_product1_12__0__q ;
wire Xd_0__inst_product1_13__0__q ;
wire Xd_0__inst_product1_14__0__q ;
wire Xd_0__inst_product1_15__0__q ;
wire Xd_0__inst_product1_10__0__q ;
wire Xd_0__inst_product1_11__0__q ;
wire Xd_0__inst_product1_8__0__q ;
wire Xd_0__inst_product1_9__0__q ;
wire Xd_0__inst_product1_6__0__q ;
wire Xd_0__inst_product1_7__0__q ;
wire Xd_0__inst_product1_4__0__q ;
wire Xd_0__inst_product1_5__0__q ;
wire Xd_0__inst_product1_2__0__q ;
wire Xd_0__inst_product1_3__0__q ;
wire Xd_0__inst_product1_0__0__q ;
wire Xd_0__inst_product1_1__0__q ;
wire Xd_0__inst_product1_12__1__q ;
wire Xd_0__inst_product1_13__1__q ;
wire Xd_0__inst_product1_14__1__q ;
wire Xd_0__inst_product1_15__1__q ;
wire Xd_0__inst_product1_10__1__q ;
wire Xd_0__inst_product1_11__1__q ;
wire Xd_0__inst_product1_8__1__q ;
wire Xd_0__inst_product1_9__1__q ;
wire Xd_0__inst_product1_6__1__q ;
wire Xd_0__inst_product1_7__1__q ;
wire Xd_0__inst_product1_4__1__q ;
wire Xd_0__inst_product1_5__1__q ;
wire Xd_0__inst_product1_2__1__q ;
wire Xd_0__inst_product1_3__1__q ;
wire Xd_0__inst_product1_0__1__q ;
wire Xd_0__inst_product1_1__1__q ;
wire Xd_0__inst_product1_12__2__q ;
wire Xd_0__inst_product1_13__2__q ;
wire Xd_0__inst_product1_14__2__q ;
wire Xd_0__inst_product1_15__2__q ;
wire Xd_0__inst_product1_10__2__q ;
wire Xd_0__inst_product1_11__2__q ;
wire Xd_0__inst_product1_8__2__q ;
wire Xd_0__inst_product1_9__2__q ;
wire Xd_0__inst_product1_6__2__q ;
wire Xd_0__inst_product1_7__2__q ;
wire Xd_0__inst_product1_4__2__q ;
wire Xd_0__inst_product1_5__2__q ;
wire Xd_0__inst_product1_2__2__q ;
wire Xd_0__inst_product1_3__2__q ;
wire Xd_0__inst_product1_0__2__q ;
wire Xd_0__inst_product1_1__2__q ;
wire Xd_0__inst_product1_12__3__q ;
wire Xd_0__inst_product1_13__3__q ;
wire Xd_0__inst_product1_14__3__q ;
wire Xd_0__inst_product1_15__3__q ;
wire Xd_0__inst_product1_10__3__q ;
wire Xd_0__inst_product1_11__3__q ;
wire Xd_0__inst_product1_8__3__q ;
wire Xd_0__inst_product1_9__3__q ;
wire Xd_0__inst_product1_6__3__q ;
wire Xd_0__inst_product1_7__3__q ;
wire Xd_0__inst_product1_4__3__q ;
wire Xd_0__inst_product1_5__3__q ;
wire Xd_0__inst_product1_2__3__q ;
wire Xd_0__inst_product1_3__3__q ;
wire Xd_0__inst_product1_0__3__q ;
wire Xd_0__inst_product1_1__3__q ;
wire Xd_0__inst_product1_12__4__q ;
wire Xd_0__inst_product1_13__4__q ;
wire Xd_0__inst_product1_14__4__q ;
wire Xd_0__inst_product1_15__4__q ;
wire Xd_0__inst_product1_10__4__q ;
wire Xd_0__inst_product1_11__4__q ;
wire Xd_0__inst_product1_8__4__q ;
wire Xd_0__inst_product1_9__4__q ;
wire Xd_0__inst_product1_6__4__q ;
wire Xd_0__inst_product1_7__4__q ;
wire Xd_0__inst_product1_4__4__q ;
wire Xd_0__inst_product1_5__4__q ;
wire Xd_0__inst_product1_2__4__q ;
wire Xd_0__inst_product1_3__4__q ;
wire Xd_0__inst_product1_0__4__q ;
wire Xd_0__inst_product1_1__4__q ;
wire Xd_0__inst_mult_12_0_q ;
wire Xd_0__inst_mult_12_1_q ;
wire Xd_0__inst_mult_13_0_q ;
wire Xd_0__inst_mult_13_1_q ;
wire Xd_0__inst_mult_14_0_q ;
wire Xd_0__inst_mult_14_1_q ;
wire Xd_0__inst_mult_15_0_q ;
wire Xd_0__inst_mult_15_1_q ;
wire Xd_0__inst_mult_10_0_q ;
wire Xd_0__inst_mult_10_1_q ;
wire Xd_0__inst_mult_11_0_q ;
wire Xd_0__inst_mult_11_1_q ;
wire Xd_0__inst_mult_8_0_q ;
wire Xd_0__inst_mult_8_1_q ;
wire Xd_0__inst_mult_9_0_q ;
wire Xd_0__inst_mult_9_1_q ;
wire Xd_0__inst_mult_6_0_q ;
wire Xd_0__inst_mult_6_1_q ;
wire Xd_0__inst_mult_7_0_q ;
wire Xd_0__inst_mult_7_1_q ;
wire Xd_0__inst_mult_4_0_q ;
wire Xd_0__inst_mult_4_1_q ;
wire Xd_0__inst_mult_5_0_q ;
wire Xd_0__inst_mult_5_1_q ;
wire Xd_0__inst_mult_2_0_q ;
wire Xd_0__inst_mult_2_1_q ;
wire Xd_0__inst_mult_3_0_q ;
wire Xd_0__inst_mult_3_1_q ;
wire Xd_0__inst_mult_0_0_q ;
wire Xd_0__inst_mult_0_1_q ;
wire Xd_0__inst_mult_1_0_q ;
wire Xd_0__inst_mult_1_1_q ;
wire Xd_0__inst_mult_12_2_q ;
wire Xd_0__inst_mult_12_3_q ;
wire Xd_0__inst_mult_13_2_q ;
wire Xd_0__inst_mult_13_3_q ;
wire Xd_0__inst_mult_14_2_q ;
wire Xd_0__inst_mult_14_3_q ;
wire Xd_0__inst_mult_15_2_q ;
wire Xd_0__inst_mult_15_3_q ;
wire Xd_0__inst_mult_10_2_q ;
wire Xd_0__inst_mult_10_3_q ;
wire Xd_0__inst_mult_11_2_q ;
wire Xd_0__inst_mult_11_3_q ;
wire Xd_0__inst_mult_8_2_q ;
wire Xd_0__inst_mult_8_3_q ;
wire Xd_0__inst_mult_9_2_q ;
wire Xd_0__inst_mult_9_3_q ;
wire Xd_0__inst_mult_6_2_q ;
wire Xd_0__inst_mult_6_3_q ;
wire Xd_0__inst_mult_7_2_q ;
wire Xd_0__inst_mult_7_3_q ;
wire Xd_0__inst_mult_4_2_q ;
wire Xd_0__inst_mult_4_3_q ;
wire Xd_0__inst_mult_5_2_q ;
wire Xd_0__inst_mult_5_3_q ;
wire Xd_0__inst_mult_2_2_q ;
wire Xd_0__inst_mult_2_3_q ;
wire Xd_0__inst_mult_3_2_q ;
wire Xd_0__inst_mult_3_3_q ;
wire Xd_0__inst_mult_0_2_q ;
wire Xd_0__inst_mult_0_3_q ;
wire Xd_0__inst_mult_1_2_q ;
wire Xd_0__inst_mult_1_3_q ;
wire Xd_0__inst_mult_12_4_q ;
wire Xd_0__inst_mult_12_5_q ;
wire Xd_0__inst_mult_13_4_q ;
wire Xd_0__inst_mult_13_5_q ;
wire Xd_0__inst_mult_14_4_q ;
wire Xd_0__inst_mult_14_5_q ;
wire Xd_0__inst_mult_15_4_q ;
wire Xd_0__inst_mult_15_5_q ;
wire Xd_0__inst_mult_10_4_q ;
wire Xd_0__inst_mult_10_5_q ;
wire Xd_0__inst_mult_11_4_q ;
wire Xd_0__inst_mult_11_5_q ;
wire Xd_0__inst_mult_8_4_q ;
wire Xd_0__inst_mult_8_5_q ;
wire Xd_0__inst_mult_9_4_q ;
wire Xd_0__inst_mult_9_5_q ;
wire Xd_0__inst_mult_6_4_q ;
wire Xd_0__inst_mult_6_5_q ;
wire Xd_0__inst_mult_7_4_q ;
wire Xd_0__inst_mult_7_5_q ;
wire Xd_0__inst_mult_4_4_q ;
wire Xd_0__inst_mult_4_5_q ;
wire Xd_0__inst_mult_5_4_q ;
wire Xd_0__inst_mult_5_5_q ;
wire Xd_0__inst_mult_2_4_q ;
wire Xd_0__inst_mult_2_5_q ;
wire Xd_0__inst_mult_3_4_q ;
wire Xd_0__inst_mult_3_5_q ;
wire Xd_0__inst_mult_0_4_q ;
wire Xd_0__inst_mult_0_5_q ;
wire Xd_0__inst_mult_1_4_q ;
wire Xd_0__inst_mult_1_5_q ;
wire Xd_0__inst_mult_12_6_q ;
wire Xd_0__inst_mult_12_7_q ;
wire Xd_0__inst_mult_13_6_q ;
wire Xd_0__inst_mult_13_7_q ;
wire Xd_0__inst_mult_14_6_q ;
wire Xd_0__inst_mult_14_7_q ;
wire Xd_0__inst_mult_15_6_q ;
wire Xd_0__inst_mult_15_7_q ;
wire Xd_0__inst_mult_10_6_q ;
wire Xd_0__inst_mult_10_7_q ;
wire Xd_0__inst_mult_11_6_q ;
wire Xd_0__inst_mult_11_7_q ;
wire Xd_0__inst_mult_8_6_q ;
wire Xd_0__inst_mult_8_7_q ;
wire Xd_0__inst_mult_9_6_q ;
wire Xd_0__inst_mult_9_7_q ;
wire Xd_0__inst_mult_6_6_q ;
wire Xd_0__inst_mult_6_7_q ;
wire Xd_0__inst_mult_7_6_q ;
wire Xd_0__inst_mult_7_7_q ;
wire Xd_0__inst_mult_4_6_q ;
wire Xd_0__inst_mult_4_7_q ;
wire Xd_0__inst_mult_5_6_q ;
wire Xd_0__inst_mult_5_7_q ;
wire Xd_0__inst_mult_2_6_q ;
wire Xd_0__inst_mult_2_7_q ;
wire Xd_0__inst_mult_3_6_q ;
wire Xd_0__inst_mult_3_7_q ;
wire Xd_0__inst_mult_0_6_q ;
wire Xd_0__inst_mult_0_7_q ;
wire Xd_0__inst_mult_1_6_q ;
wire Xd_0__inst_mult_1_7_q ;
wire Xd_0__inst_mult_12_8_q ;
wire Xd_0__inst_mult_12_9_q ;
wire Xd_0__inst_mult_13_8_q ;
wire Xd_0__inst_mult_13_9_q ;
wire Xd_0__inst_mult_14_8_q ;
wire Xd_0__inst_mult_14_9_q ;
wire Xd_0__inst_mult_15_8_q ;
wire Xd_0__inst_mult_15_9_q ;
wire Xd_0__inst_mult_10_8_q ;
wire Xd_0__inst_mult_10_9_q ;
wire Xd_0__inst_mult_11_8_q ;
wire Xd_0__inst_mult_11_9_q ;
wire Xd_0__inst_mult_8_8_q ;
wire Xd_0__inst_mult_8_9_q ;
wire Xd_0__inst_mult_9_8_q ;
wire Xd_0__inst_mult_9_9_q ;
wire Xd_0__inst_mult_6_8_q ;
wire Xd_0__inst_mult_6_9_q ;
wire Xd_0__inst_mult_7_8_q ;
wire Xd_0__inst_mult_7_9_q ;
wire Xd_0__inst_mult_4_8_q ;
wire Xd_0__inst_mult_4_9_q ;
wire Xd_0__inst_mult_5_8_q ;
wire Xd_0__inst_mult_5_9_q ;
wire Xd_0__inst_mult_2_8_q ;
wire Xd_0__inst_mult_2_9_q ;
wire Xd_0__inst_mult_3_8_q ;
wire Xd_0__inst_mult_3_9_q ;
wire Xd_0__inst_mult_0_8_q ;
wire Xd_0__inst_mult_0_9_q ;
wire Xd_0__inst_mult_1_8_q ;
wire Xd_0__inst_mult_1_9_q ;
wire Xd_0__inst_mult_12_10_q ;
wire Xd_0__inst_mult_12_11_q ;
wire Xd_0__inst_mult_13_10_q ;
wire Xd_0__inst_mult_13_11_q ;
wire Xd_0__inst_mult_14_10_q ;
wire Xd_0__inst_mult_14_11_q ;
wire Xd_0__inst_mult_15_10_q ;
wire Xd_0__inst_mult_15_11_q ;
wire Xd_0__inst_mult_10_10_q ;
wire Xd_0__inst_mult_10_11_q ;
wire Xd_0__inst_mult_11_10_q ;
wire Xd_0__inst_mult_11_11_q ;
wire Xd_0__inst_mult_8_10_q ;
wire Xd_0__inst_mult_8_11_q ;
wire Xd_0__inst_mult_9_10_q ;
wire Xd_0__inst_mult_9_11_q ;
wire Xd_0__inst_mult_6_10_q ;
wire Xd_0__inst_mult_6_11_q ;
wire Xd_0__inst_mult_7_10_q ;
wire Xd_0__inst_mult_7_11_q ;
wire Xd_0__inst_mult_4_10_q ;
wire Xd_0__inst_mult_4_11_q ;
wire Xd_0__inst_mult_5_10_q ;
wire Xd_0__inst_mult_5_11_q ;
wire Xd_0__inst_mult_2_10_q ;
wire Xd_0__inst_mult_2_11_q ;
wire Xd_0__inst_mult_3_10_q ;
wire Xd_0__inst_mult_3_11_q ;
wire Xd_0__inst_mult_0_10_q ;
wire Xd_0__inst_mult_0_11_q ;
wire Xd_0__inst_mult_1_10_q ;
wire Xd_0__inst_mult_1_11_q ;
wire Xd_0__inst_mult_12_12_q ;
wire Xd_0__inst_mult_12_13_q ;
wire Xd_0__inst_mult_13_12_q ;
wire Xd_0__inst_mult_13_13_q ;
wire Xd_0__inst_mult_14_12_q ;
wire Xd_0__inst_mult_14_13_q ;
wire Xd_0__inst_mult_15_12_q ;
wire Xd_0__inst_mult_15_13_q ;
wire Xd_0__inst_mult_10_12_q ;
wire Xd_0__inst_mult_10_13_q ;
wire Xd_0__inst_mult_11_12_q ;
wire Xd_0__inst_mult_11_13_q ;
wire Xd_0__inst_mult_8_12_q ;
wire Xd_0__inst_mult_8_13_q ;
wire Xd_0__inst_mult_9_12_q ;
wire Xd_0__inst_mult_9_13_q ;
wire Xd_0__inst_mult_6_12_q ;
wire Xd_0__inst_mult_6_13_q ;
wire Xd_0__inst_mult_7_12_q ;
wire Xd_0__inst_mult_7_13_q ;
wire Xd_0__inst_mult_4_12_q ;
wire Xd_0__inst_mult_4_13_q ;
wire Xd_0__inst_mult_5_12_q ;
wire Xd_0__inst_mult_5_13_q ;
wire Xd_0__inst_mult_2_12_q ;
wire Xd_0__inst_mult_2_13_q ;
wire Xd_0__inst_mult_3_12_q ;
wire Xd_0__inst_mult_3_13_q ;
wire Xd_0__inst_mult_0_12_q ;
wire Xd_0__inst_mult_0_13_q ;
wire Xd_0__inst_mult_1_12_q ;
wire Xd_0__inst_mult_1_13_q ;
wire Xd_0__inst_mult_12_14_q ;
wire Xd_0__inst_mult_12_15_q ;
wire Xd_0__inst_mult_13_14_q ;
wire Xd_0__inst_mult_13_15_q ;
wire Xd_0__inst_mult_14_14_q ;
wire Xd_0__inst_mult_14_15_q ;
wire Xd_0__inst_mult_15_14_q ;
wire Xd_0__inst_mult_15_15_q ;
wire Xd_0__inst_mult_10_14_q ;
wire Xd_0__inst_mult_10_15_q ;
wire Xd_0__inst_mult_11_14_q ;
wire Xd_0__inst_mult_11_15_q ;
wire Xd_0__inst_mult_8_14_q ;
wire Xd_0__inst_mult_8_15_q ;
wire Xd_0__inst_mult_9_14_q ;
wire Xd_0__inst_mult_9_15_q ;
wire Xd_0__inst_mult_6_14_q ;
wire Xd_0__inst_mult_6_15_q ;
wire Xd_0__inst_mult_7_14_q ;
wire Xd_0__inst_mult_7_15_q ;
wire Xd_0__inst_mult_4_14_q ;
wire Xd_0__inst_mult_4_15_q ;
wire Xd_0__inst_mult_5_14_q ;
wire Xd_0__inst_mult_5_15_q ;
wire Xd_0__inst_mult_2_14_q ;
wire Xd_0__inst_mult_2_15_q ;
wire Xd_0__inst_mult_3_14_q ;
wire Xd_0__inst_mult_3_15_q ;
wire Xd_0__inst_mult_0_14_q ;
wire Xd_0__inst_mult_0_15_q ;
wire Xd_0__inst_mult_1_14_q ;
wire Xd_0__inst_mult_1_15_q ;
wire Xd_0__inst_mult_12_16_q ;
wire Xd_0__inst_mult_12_17_q ;
wire Xd_0__inst_mult_13_16_q ;
wire Xd_0__inst_mult_13_17_q ;
wire Xd_0__inst_mult_14_16_q ;
wire Xd_0__inst_mult_14_17_q ;
wire Xd_0__inst_mult_15_16_q ;
wire Xd_0__inst_mult_15_17_q ;
wire Xd_0__inst_mult_10_16_q ;
wire Xd_0__inst_mult_10_17_q ;
wire Xd_0__inst_mult_11_16_q ;
wire Xd_0__inst_mult_11_17_q ;
wire Xd_0__inst_mult_8_16_q ;
wire Xd_0__inst_mult_8_17_q ;
wire Xd_0__inst_mult_9_16_q ;
wire Xd_0__inst_mult_9_17_q ;
wire Xd_0__inst_mult_6_16_q ;
wire Xd_0__inst_mult_6_17_q ;
wire Xd_0__inst_mult_7_16_q ;
wire Xd_0__inst_mult_7_17_q ;
wire Xd_0__inst_mult_4_16_q ;
wire Xd_0__inst_mult_4_17_q ;
wire Xd_0__inst_mult_5_16_q ;
wire Xd_0__inst_mult_5_17_q ;
wire Xd_0__inst_mult_2_16_q ;
wire Xd_0__inst_mult_2_17_q ;
wire Xd_0__inst_mult_3_16_q ;
wire Xd_0__inst_mult_3_17_q ;
wire Xd_0__inst_mult_0_16_q ;
wire Xd_0__inst_mult_0_17_q ;
wire Xd_0__inst_mult_1_16_q ;
wire Xd_0__inst_mult_1_17_q ;
wire Xd_0__inst_mult_12_18_q ;
wire Xd_0__inst_mult_12_19_q ;
wire Xd_0__inst_mult_13_18_q ;
wire Xd_0__inst_mult_13_19_q ;
wire Xd_0__inst_mult_14_18_q ;
wire Xd_0__inst_mult_14_19_q ;
wire Xd_0__inst_mult_15_18_q ;
wire Xd_0__inst_mult_15_19_q ;
wire Xd_0__inst_mult_10_18_q ;
wire Xd_0__inst_mult_10_19_q ;
wire Xd_0__inst_mult_11_18_q ;
wire Xd_0__inst_mult_11_19_q ;
wire Xd_0__inst_mult_8_18_q ;
wire Xd_0__inst_mult_8_19_q ;
wire Xd_0__inst_mult_9_18_q ;
wire Xd_0__inst_mult_9_19_q ;
wire Xd_0__inst_mult_6_18_q ;
wire Xd_0__inst_mult_6_19_q ;
wire Xd_0__inst_mult_7_18_q ;
wire Xd_0__inst_mult_7_19_q ;
wire Xd_0__inst_mult_4_18_q ;
wire Xd_0__inst_mult_4_19_q ;
wire Xd_0__inst_mult_5_18_q ;
wire Xd_0__inst_mult_5_19_q ;
wire Xd_0__inst_mult_2_18_q ;
wire Xd_0__inst_mult_2_19_q ;
wire Xd_0__inst_mult_3_18_q ;
wire Xd_0__inst_mult_3_19_q ;
wire Xd_0__inst_mult_0_18_q ;
wire Xd_0__inst_mult_0_19_q ;
wire Xd_0__inst_mult_1_18_q ;
wire Xd_0__inst_mult_1_19_q ;
wire Xd_0__inst_mult_12_20_q ;
wire Xd_0__inst_mult_12_21_q ;
wire Xd_0__inst_mult_12_22_q ;
wire Xd_0__inst_mult_12_23_q ;
wire Xd_0__inst_mult_13_20_q ;
wire Xd_0__inst_mult_13_21_q ;
wire Xd_0__inst_mult_13_22_q ;
wire Xd_0__inst_mult_13_23_q ;
wire Xd_0__inst_mult_14_20_q ;
wire Xd_0__inst_mult_14_21_q ;
wire Xd_0__inst_mult_14_22_q ;
wire Xd_0__inst_mult_14_23_q ;
wire Xd_0__inst_mult_15_20_q ;
wire Xd_0__inst_mult_15_21_q ;
wire Xd_0__inst_mult_15_22_q ;
wire Xd_0__inst_mult_15_23_q ;
wire Xd_0__inst_mult_10_20_q ;
wire Xd_0__inst_mult_10_21_q ;
wire Xd_0__inst_mult_10_22_q ;
wire Xd_0__inst_mult_10_23_q ;
wire Xd_0__inst_mult_11_20_q ;
wire Xd_0__inst_mult_11_21_q ;
wire Xd_0__inst_mult_11_22_q ;
wire Xd_0__inst_mult_11_23_q ;
wire Xd_0__inst_mult_8_20_q ;
wire Xd_0__inst_mult_8_21_q ;
wire Xd_0__inst_mult_8_22_q ;
wire Xd_0__inst_mult_8_23_q ;
wire Xd_0__inst_mult_9_20_q ;
wire Xd_0__inst_mult_9_21_q ;
wire Xd_0__inst_mult_9_22_q ;
wire Xd_0__inst_mult_9_23_q ;
wire Xd_0__inst_mult_6_20_q ;
wire Xd_0__inst_mult_6_21_q ;
wire Xd_0__inst_mult_6_22_q ;
wire Xd_0__inst_mult_6_23_q ;
wire Xd_0__inst_mult_7_20_q ;
wire Xd_0__inst_mult_7_21_q ;
wire Xd_0__inst_mult_7_22_q ;
wire Xd_0__inst_mult_7_23_q ;
wire Xd_0__inst_mult_4_20_q ;
wire Xd_0__inst_mult_4_21_q ;
wire Xd_0__inst_mult_4_22_q ;
wire Xd_0__inst_mult_4_23_q ;
wire Xd_0__inst_mult_5_20_q ;
wire Xd_0__inst_mult_5_21_q ;
wire Xd_0__inst_mult_5_22_q ;
wire Xd_0__inst_mult_5_23_q ;
wire Xd_0__inst_mult_2_20_q ;
wire Xd_0__inst_mult_2_21_q ;
wire Xd_0__inst_mult_2_22_q ;
wire Xd_0__inst_mult_2_23_q ;
wire Xd_0__inst_mult_3_20_q ;
wire Xd_0__inst_mult_3_21_q ;
wire Xd_0__inst_mult_3_22_q ;
wire Xd_0__inst_mult_3_23_q ;
wire Xd_0__inst_mult_0_20_q ;
wire Xd_0__inst_mult_0_21_q ;
wire Xd_0__inst_mult_0_22_q ;
wire Xd_0__inst_mult_0_23_q ;
wire Xd_0__inst_mult_1_20_q ;
wire Xd_0__inst_mult_1_21_q ;
wire Xd_0__inst_mult_1_22_q ;
wire Xd_0__inst_mult_1_23_q ;
wire Xd_0__inst_mult_12_24_q ;
wire Xd_0__inst_mult_12_25_q ;
wire Xd_0__inst_mult_13_24_q ;
wire Xd_0__inst_mult_13_25_q ;
wire Xd_0__inst_mult_14_24_q ;
wire Xd_0__inst_mult_14_25_q ;
wire Xd_0__inst_mult_15_24_q ;
wire Xd_0__inst_mult_15_25_q ;
wire Xd_0__inst_mult_10_24_q ;
wire Xd_0__inst_mult_10_25_q ;
wire Xd_0__inst_mult_11_24_q ;
wire Xd_0__inst_mult_11_25_q ;
wire Xd_0__inst_mult_8_24_q ;
wire Xd_0__inst_mult_8_25_q ;
wire Xd_0__inst_mult_9_24_q ;
wire Xd_0__inst_mult_9_25_q ;
wire Xd_0__inst_mult_6_24_q ;
wire Xd_0__inst_mult_6_25_q ;
wire Xd_0__inst_mult_7_24_q ;
wire Xd_0__inst_mult_7_25_q ;
wire Xd_0__inst_mult_4_24_q ;
wire Xd_0__inst_mult_4_25_q ;
wire Xd_0__inst_mult_5_24_q ;
wire Xd_0__inst_mult_5_25_q ;
wire Xd_0__inst_mult_2_24_q ;
wire Xd_0__inst_mult_2_25_q ;
wire Xd_0__inst_mult_3_24_q ;
wire Xd_0__inst_mult_3_25_q ;
wire Xd_0__inst_mult_0_24_q ;
wire Xd_0__inst_mult_0_25_q ;
wire Xd_0__inst_mult_1_24_q ;
wire Xd_0__inst_mult_1_25_q ;
wire Xd_0__inst_mult_12_26_q ;
wire Xd_0__inst_mult_12_27_q ;
wire Xd_0__inst_mult_13_26_q ;
wire Xd_0__inst_mult_13_27_q ;
wire Xd_0__inst_mult_14_26_q ;
wire Xd_0__inst_mult_14_27_q ;
wire Xd_0__inst_mult_15_26_q ;
wire Xd_0__inst_mult_15_27_q ;
wire Xd_0__inst_mult_10_26_q ;
wire Xd_0__inst_mult_10_27_q ;
wire Xd_0__inst_mult_11_26_q ;
wire Xd_0__inst_mult_11_27_q ;
wire Xd_0__inst_mult_8_26_q ;
wire Xd_0__inst_mult_8_27_q ;
wire Xd_0__inst_mult_9_26_q ;
wire Xd_0__inst_mult_9_27_q ;
wire Xd_0__inst_mult_6_26_q ;
wire Xd_0__inst_mult_6_27_q ;
wire Xd_0__inst_mult_7_26_q ;
wire Xd_0__inst_mult_7_27_q ;
wire Xd_0__inst_mult_4_26_q ;
wire Xd_0__inst_mult_4_27_q ;
wire Xd_0__inst_mult_5_26_q ;
wire Xd_0__inst_mult_5_27_q ;
wire Xd_0__inst_mult_2_26_q ;
wire Xd_0__inst_mult_2_27_q ;
wire Xd_0__inst_mult_3_26_q ;
wire Xd_0__inst_mult_3_27_q ;
wire Xd_0__inst_mult_0_26_q ;
wire Xd_0__inst_mult_0_27_q ;
wire Xd_0__inst_mult_1_26_q ;
wire Xd_0__inst_mult_1_27_q ;
wire Xd_0__inst_mult_12_28_q ;
wire Xd_0__inst_mult_12_29_q ;
wire Xd_0__inst_mult_13_28_q ;
wire Xd_0__inst_mult_13_29_q ;
wire Xd_0__inst_mult_14_28_q ;
wire Xd_0__inst_mult_14_29_q ;
wire Xd_0__inst_mult_15_28_q ;
wire Xd_0__inst_mult_15_29_q ;
wire Xd_0__inst_mult_10_28_q ;
wire Xd_0__inst_mult_10_29_q ;
wire Xd_0__inst_mult_11_28_q ;
wire Xd_0__inst_mult_11_29_q ;
wire Xd_0__inst_mult_8_28_q ;
wire Xd_0__inst_mult_8_29_q ;
wire Xd_0__inst_mult_9_28_q ;
wire Xd_0__inst_mult_9_29_q ;
wire Xd_0__inst_mult_6_28_q ;
wire Xd_0__inst_mult_6_29_q ;
wire Xd_0__inst_mult_7_28_q ;
wire Xd_0__inst_mult_7_29_q ;
wire Xd_0__inst_mult_4_28_q ;
wire Xd_0__inst_mult_4_29_q ;
wire Xd_0__inst_mult_5_28_q ;
wire Xd_0__inst_mult_5_29_q ;
wire Xd_0__inst_mult_2_28_q ;
wire Xd_0__inst_mult_2_29_q ;
wire Xd_0__inst_mult_3_28_q ;
wire Xd_0__inst_mult_3_29_q ;
wire Xd_0__inst_mult_0_28_q ;
wire Xd_0__inst_mult_0_29_q ;
wire Xd_0__inst_mult_1_28_q ;
wire Xd_0__inst_mult_1_29_q ;
wire Xd_0__inst_mult_12_30_q ;
wire Xd_0__inst_mult_12_31_q ;
wire Xd_0__inst_mult_13_30_q ;
wire Xd_0__inst_mult_13_31_q ;
wire Xd_0__inst_mult_14_30_q ;
wire Xd_0__inst_mult_14_31_q ;
wire Xd_0__inst_mult_15_30_q ;
wire Xd_0__inst_mult_15_31_q ;
wire Xd_0__inst_mult_10_30_q ;
wire Xd_0__inst_mult_10_31_q ;
wire Xd_0__inst_mult_11_30_q ;
wire Xd_0__inst_mult_11_31_q ;
wire Xd_0__inst_mult_8_30_q ;
wire Xd_0__inst_mult_8_31_q ;
wire Xd_0__inst_mult_9_30_q ;
wire Xd_0__inst_mult_9_31_q ;
wire Xd_0__inst_mult_6_30_q ;
wire Xd_0__inst_mult_6_31_q ;
wire Xd_0__inst_mult_7_30_q ;
wire Xd_0__inst_mult_7_31_q ;
wire Xd_0__inst_mult_4_30_q ;
wire Xd_0__inst_mult_4_31_q ;
wire Xd_0__inst_mult_5_30_q ;
wire Xd_0__inst_mult_5_31_q ;
wire Xd_0__inst_mult_2_30_q ;
wire Xd_0__inst_mult_2_31_q ;
wire Xd_0__inst_mult_3_30_q ;
wire Xd_0__inst_mult_3_31_q ;
wire Xd_0__inst_mult_0_30_q ;
wire Xd_0__inst_mult_0_31_q ;
wire Xd_0__inst_mult_1_30_q ;
wire Xd_0__inst_mult_1_31_q ;
wire Xd_0__inst_mult_12_32_q ;
wire Xd_0__inst_mult_12_33_q ;
wire Xd_0__inst_mult_13_32_q ;
wire Xd_0__inst_mult_13_33_q ;
wire Xd_0__inst_mult_14_32_q ;
wire Xd_0__inst_mult_14_33_q ;
wire Xd_0__inst_mult_15_32_q ;
wire Xd_0__inst_mult_15_33_q ;
wire Xd_0__inst_mult_10_32_q ;
wire Xd_0__inst_mult_10_33_q ;
wire Xd_0__inst_mult_11_32_q ;
wire Xd_0__inst_mult_11_33_q ;
wire Xd_0__inst_mult_8_32_q ;
wire Xd_0__inst_mult_8_33_q ;
wire Xd_0__inst_mult_9_32_q ;
wire Xd_0__inst_mult_9_33_q ;
wire Xd_0__inst_mult_6_32_q ;
wire Xd_0__inst_mult_6_33_q ;
wire Xd_0__inst_mult_7_32_q ;
wire Xd_0__inst_mult_7_33_q ;
wire Xd_0__inst_mult_4_32_q ;
wire Xd_0__inst_mult_4_33_q ;
wire Xd_0__inst_mult_5_32_q ;
wire Xd_0__inst_mult_5_33_q ;
wire Xd_0__inst_mult_2_32_q ;
wire Xd_0__inst_mult_2_33_q ;
wire Xd_0__inst_mult_3_32_q ;
wire Xd_0__inst_mult_3_33_q ;
wire Xd_0__inst_mult_0_32_q ;
wire Xd_0__inst_mult_0_33_q ;
wire Xd_0__inst_mult_1_32_q ;
wire Xd_0__inst_mult_1_33_q ;
wire [0:15] Xd_0__inst_sign1 ;
wire [23:0] Xd_0__inst_a1_4__adder1_inst_dout ;
wire [0:15] Xd_0__inst_sign ;
wire [23:0] Xd_0__inst_a1_5__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_7__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_6__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_3__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_2__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_1__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_0__adder1_inst_dout ;
wire [26:0] Xd_0__inst_inst_inst_dout ;


twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_1 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_1_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q  $ (Xd_0__inst_inst_first_level_0__0__q )) ) + ( Xd_0__inst_mult_4_175  ) + ( Xd_0__inst_mult_4_174  ))
// Xd_0__inst_inst_inst_rtl_2  = CARRY(( !Xd_0__inst_inst_first_level_2__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q  $ (Xd_0__inst_inst_first_level_0__0__q )) ) + ( Xd_0__inst_mult_4_175  ) + ( Xd_0__inst_mult_4_174  ))
// Xd_0__inst_inst_inst_rtl_3  = SHARE((!Xd_0__inst_inst_first_level_2__0__q  & (Xd_0__inst_inst_first_level_1__0__q  & Xd_0__inst_inst_first_level_0__0__q )) # (Xd_0__inst_inst_first_level_2__0__q  & ((Xd_0__inst_inst_first_level_0__0__q ) # 
// (Xd_0__inst_inst_first_level_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__0__q ),
	.datac(!Xd_0__inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_174 ),
	.sharein(Xd_0__inst_mult_4_175 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_1_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_2 ),
	.shareout(Xd_0__inst_inst_inst_rtl_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_5 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_5_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q  $ (Xd_0__inst_inst_first_level_0__1__q )) ) + ( Xd_0__inst_inst_inst_rtl_3  ) + ( Xd_0__inst_inst_inst_rtl_2  ))
// Xd_0__inst_inst_inst_rtl_6  = CARRY(( !Xd_0__inst_inst_first_level_2__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q  $ (Xd_0__inst_inst_first_level_0__1__q )) ) + ( Xd_0__inst_inst_inst_rtl_3  ) + ( Xd_0__inst_inst_inst_rtl_2  ))
// Xd_0__inst_inst_inst_rtl_7  = SHARE((!Xd_0__inst_inst_first_level_2__1__q  & (Xd_0__inst_inst_first_level_1__1__q  & Xd_0__inst_inst_first_level_0__1__q )) # (Xd_0__inst_inst_first_level_2__1__q  & ((Xd_0__inst_inst_first_level_0__1__q ) # 
// (Xd_0__inst_inst_first_level_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__1__q ),
	.datac(!Xd_0__inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_2 ),
	.sharein(Xd_0__inst_inst_inst_rtl_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_5_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_6 ),
	.shareout(Xd_0__inst_inst_inst_rtl_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_9 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_9_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q  $ (Xd_0__inst_inst_first_level_0__2__q )) ) + ( Xd_0__inst_inst_inst_rtl_7  ) + ( Xd_0__inst_inst_inst_rtl_6  ))
// Xd_0__inst_inst_inst_rtl_10  = CARRY(( !Xd_0__inst_inst_first_level_2__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q  $ (Xd_0__inst_inst_first_level_0__2__q )) ) + ( Xd_0__inst_inst_inst_rtl_7  ) + ( Xd_0__inst_inst_inst_rtl_6  ))
// Xd_0__inst_inst_inst_rtl_11  = SHARE((!Xd_0__inst_inst_first_level_2__2__q  & (Xd_0__inst_inst_first_level_1__2__q  & Xd_0__inst_inst_first_level_0__2__q )) # (Xd_0__inst_inst_first_level_2__2__q  & ((Xd_0__inst_inst_first_level_0__2__q ) # 
// (Xd_0__inst_inst_first_level_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__2__q ),
	.datac(!Xd_0__inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_6 ),
	.sharein(Xd_0__inst_inst_inst_rtl_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_9_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_10 ),
	.shareout(Xd_0__inst_inst_inst_rtl_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_13 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_13_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q  $ (Xd_0__inst_inst_first_level_0__3__q )) ) + ( Xd_0__inst_inst_inst_rtl_11  ) + ( Xd_0__inst_inst_inst_rtl_10  ))
// Xd_0__inst_inst_inst_rtl_14  = CARRY(( !Xd_0__inst_inst_first_level_2__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q  $ (Xd_0__inst_inst_first_level_0__3__q )) ) + ( Xd_0__inst_inst_inst_rtl_11  ) + ( Xd_0__inst_inst_inst_rtl_10  ))
// Xd_0__inst_inst_inst_rtl_15  = SHARE((!Xd_0__inst_inst_first_level_2__3__q  & (Xd_0__inst_inst_first_level_1__3__q  & Xd_0__inst_inst_first_level_0__3__q )) # (Xd_0__inst_inst_first_level_2__3__q  & ((Xd_0__inst_inst_first_level_0__3__q ) # 
// (Xd_0__inst_inst_first_level_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__3__q ),
	.datac(!Xd_0__inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_10 ),
	.sharein(Xd_0__inst_inst_inst_rtl_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_13_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_14 ),
	.shareout(Xd_0__inst_inst_inst_rtl_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_17 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_17_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q  $ (Xd_0__inst_inst_first_level_0__4__q )) ) + ( Xd_0__inst_inst_inst_rtl_15  ) + ( Xd_0__inst_inst_inst_rtl_14  ))
// Xd_0__inst_inst_inst_rtl_18  = CARRY(( !Xd_0__inst_inst_first_level_2__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q  $ (Xd_0__inst_inst_first_level_0__4__q )) ) + ( Xd_0__inst_inst_inst_rtl_15  ) + ( Xd_0__inst_inst_inst_rtl_14  ))
// Xd_0__inst_inst_inst_rtl_19  = SHARE((!Xd_0__inst_inst_first_level_2__4__q  & (Xd_0__inst_inst_first_level_1__4__q  & Xd_0__inst_inst_first_level_0__4__q )) # (Xd_0__inst_inst_first_level_2__4__q  & ((Xd_0__inst_inst_first_level_0__4__q ) # 
// (Xd_0__inst_inst_first_level_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__4__q ),
	.datac(!Xd_0__inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_14 ),
	.sharein(Xd_0__inst_inst_inst_rtl_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_17_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_18 ),
	.shareout(Xd_0__inst_inst_inst_rtl_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_21 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_21_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q  $ (Xd_0__inst_inst_first_level_0__5__q )) ) + ( Xd_0__inst_inst_inst_rtl_19  ) + ( Xd_0__inst_inst_inst_rtl_18  ))
// Xd_0__inst_inst_inst_rtl_22  = CARRY(( !Xd_0__inst_inst_first_level_2__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q  $ (Xd_0__inst_inst_first_level_0__5__q )) ) + ( Xd_0__inst_inst_inst_rtl_19  ) + ( Xd_0__inst_inst_inst_rtl_18  ))
// Xd_0__inst_inst_inst_rtl_23  = SHARE((!Xd_0__inst_inst_first_level_2__5__q  & (Xd_0__inst_inst_first_level_1__5__q  & Xd_0__inst_inst_first_level_0__5__q )) # (Xd_0__inst_inst_first_level_2__5__q  & ((Xd_0__inst_inst_first_level_0__5__q ) # 
// (Xd_0__inst_inst_first_level_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__5__q ),
	.datac(!Xd_0__inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_18 ),
	.sharein(Xd_0__inst_inst_inst_rtl_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_21_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_22 ),
	.shareout(Xd_0__inst_inst_inst_rtl_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_25 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_25_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q  $ (Xd_0__inst_inst_first_level_0__6__q )) ) + ( Xd_0__inst_inst_inst_rtl_23  ) + ( Xd_0__inst_inst_inst_rtl_22  ))
// Xd_0__inst_inst_inst_rtl_26  = CARRY(( !Xd_0__inst_inst_first_level_2__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q  $ (Xd_0__inst_inst_first_level_0__6__q )) ) + ( Xd_0__inst_inst_inst_rtl_23  ) + ( Xd_0__inst_inst_inst_rtl_22  ))
// Xd_0__inst_inst_inst_rtl_27  = SHARE((!Xd_0__inst_inst_first_level_2__6__q  & (Xd_0__inst_inst_first_level_1__6__q  & Xd_0__inst_inst_first_level_0__6__q )) # (Xd_0__inst_inst_first_level_2__6__q  & ((Xd_0__inst_inst_first_level_0__6__q ) # 
// (Xd_0__inst_inst_first_level_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__6__q ),
	.datac(!Xd_0__inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_22 ),
	.sharein(Xd_0__inst_inst_inst_rtl_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_25_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_26 ),
	.shareout(Xd_0__inst_inst_inst_rtl_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_29 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_29_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q  $ (Xd_0__inst_inst_first_level_0__7__q )) ) + ( Xd_0__inst_inst_inst_rtl_27  ) + ( Xd_0__inst_inst_inst_rtl_26  ))
// Xd_0__inst_inst_inst_rtl_30  = CARRY(( !Xd_0__inst_inst_first_level_2__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q  $ (Xd_0__inst_inst_first_level_0__7__q )) ) + ( Xd_0__inst_inst_inst_rtl_27  ) + ( Xd_0__inst_inst_inst_rtl_26  ))
// Xd_0__inst_inst_inst_rtl_31  = SHARE((!Xd_0__inst_inst_first_level_2__7__q  & (Xd_0__inst_inst_first_level_1__7__q  & Xd_0__inst_inst_first_level_0__7__q )) # (Xd_0__inst_inst_first_level_2__7__q  & ((Xd_0__inst_inst_first_level_0__7__q ) # 
// (Xd_0__inst_inst_first_level_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__7__q ),
	.datac(!Xd_0__inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_26 ),
	.sharein(Xd_0__inst_inst_inst_rtl_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_29_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_30 ),
	.shareout(Xd_0__inst_inst_inst_rtl_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_33 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_33_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q  $ (Xd_0__inst_inst_first_level_0__8__q )) ) + ( Xd_0__inst_inst_inst_rtl_31  ) + ( Xd_0__inst_inst_inst_rtl_30  ))
// Xd_0__inst_inst_inst_rtl_34  = CARRY(( !Xd_0__inst_inst_first_level_2__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q  $ (Xd_0__inst_inst_first_level_0__8__q )) ) + ( Xd_0__inst_inst_inst_rtl_31  ) + ( Xd_0__inst_inst_inst_rtl_30  ))
// Xd_0__inst_inst_inst_rtl_35  = SHARE((!Xd_0__inst_inst_first_level_2__8__q  & (Xd_0__inst_inst_first_level_1__8__q  & Xd_0__inst_inst_first_level_0__8__q )) # (Xd_0__inst_inst_first_level_2__8__q  & ((Xd_0__inst_inst_first_level_0__8__q ) # 
// (Xd_0__inst_inst_first_level_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__8__q ),
	.datac(!Xd_0__inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_30 ),
	.sharein(Xd_0__inst_inst_inst_rtl_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_33_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_34 ),
	.shareout(Xd_0__inst_inst_inst_rtl_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_37 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_37_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q  $ (Xd_0__inst_inst_first_level_0__9__q )) ) + ( Xd_0__inst_inst_inst_rtl_35  ) + ( Xd_0__inst_inst_inst_rtl_34  ))
// Xd_0__inst_inst_inst_rtl_38  = CARRY(( !Xd_0__inst_inst_first_level_2__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q  $ (Xd_0__inst_inst_first_level_0__9__q )) ) + ( Xd_0__inst_inst_inst_rtl_35  ) + ( Xd_0__inst_inst_inst_rtl_34  ))
// Xd_0__inst_inst_inst_rtl_39  = SHARE((!Xd_0__inst_inst_first_level_2__9__q  & (Xd_0__inst_inst_first_level_1__9__q  & Xd_0__inst_inst_first_level_0__9__q )) # (Xd_0__inst_inst_first_level_2__9__q  & ((Xd_0__inst_inst_first_level_0__9__q ) # 
// (Xd_0__inst_inst_first_level_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__9__q ),
	.datac(!Xd_0__inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_34 ),
	.sharein(Xd_0__inst_inst_inst_rtl_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_37_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_38 ),
	.shareout(Xd_0__inst_inst_inst_rtl_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_41 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_41_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q  $ (Xd_0__inst_inst_first_level_0__10__q )) ) + ( Xd_0__inst_inst_inst_rtl_39  ) + ( Xd_0__inst_inst_inst_rtl_38  ))
// Xd_0__inst_inst_inst_rtl_42  = CARRY(( !Xd_0__inst_inst_first_level_2__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q  $ (Xd_0__inst_inst_first_level_0__10__q )) ) + ( Xd_0__inst_inst_inst_rtl_39  ) + ( Xd_0__inst_inst_inst_rtl_38  ))
// Xd_0__inst_inst_inst_rtl_43  = SHARE((!Xd_0__inst_inst_first_level_2__10__q  & (Xd_0__inst_inst_first_level_1__10__q  & Xd_0__inst_inst_first_level_0__10__q )) # (Xd_0__inst_inst_first_level_2__10__q  & ((Xd_0__inst_inst_first_level_0__10__q ) # 
// (Xd_0__inst_inst_first_level_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__10__q ),
	.datac(!Xd_0__inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_38 ),
	.sharein(Xd_0__inst_inst_inst_rtl_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_41_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_42 ),
	.shareout(Xd_0__inst_inst_inst_rtl_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_45 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_45_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q  $ (Xd_0__inst_inst_first_level_0__11__q )) ) + ( Xd_0__inst_inst_inst_rtl_43  ) + ( Xd_0__inst_inst_inst_rtl_42  ))
// Xd_0__inst_inst_inst_rtl_46  = CARRY(( !Xd_0__inst_inst_first_level_2__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q  $ (Xd_0__inst_inst_first_level_0__11__q )) ) + ( Xd_0__inst_inst_inst_rtl_43  ) + ( Xd_0__inst_inst_inst_rtl_42  ))
// Xd_0__inst_inst_inst_rtl_47  = SHARE((!Xd_0__inst_inst_first_level_2__11__q  & (Xd_0__inst_inst_first_level_1__11__q  & Xd_0__inst_inst_first_level_0__11__q )) # (Xd_0__inst_inst_first_level_2__11__q  & ((Xd_0__inst_inst_first_level_0__11__q ) # 
// (Xd_0__inst_inst_first_level_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__11__q ),
	.datac(!Xd_0__inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_42 ),
	.sharein(Xd_0__inst_inst_inst_rtl_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_45_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_46 ),
	.shareout(Xd_0__inst_inst_inst_rtl_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_49 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_49_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q  $ (Xd_0__inst_inst_first_level_0__12__q )) ) + ( Xd_0__inst_inst_inst_rtl_47  ) + ( Xd_0__inst_inst_inst_rtl_46  ))
// Xd_0__inst_inst_inst_rtl_50  = CARRY(( !Xd_0__inst_inst_first_level_2__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q  $ (Xd_0__inst_inst_first_level_0__12__q )) ) + ( Xd_0__inst_inst_inst_rtl_47  ) + ( Xd_0__inst_inst_inst_rtl_46  ))
// Xd_0__inst_inst_inst_rtl_51  = SHARE((!Xd_0__inst_inst_first_level_2__12__q  & (Xd_0__inst_inst_first_level_1__12__q  & Xd_0__inst_inst_first_level_0__12__q )) # (Xd_0__inst_inst_first_level_2__12__q  & ((Xd_0__inst_inst_first_level_0__12__q ) # 
// (Xd_0__inst_inst_first_level_1__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__12__q ),
	.datac(!Xd_0__inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_46 ),
	.sharein(Xd_0__inst_inst_inst_rtl_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_49_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_50 ),
	.shareout(Xd_0__inst_inst_inst_rtl_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_53 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_53_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_rtl_51  ) + ( Xd_0__inst_inst_inst_rtl_50  ))
// Xd_0__inst_inst_inst_rtl_54  = CARRY(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_rtl_51  ) + ( Xd_0__inst_inst_inst_rtl_50  ))
// Xd_0__inst_inst_inst_rtl_55  = SHARE((!Xd_0__inst_inst_first_level_2__13__q  & (Xd_0__inst_inst_first_level_1__13__q  & Xd_0__inst_inst_first_level_0__13__q )) # (Xd_0__inst_inst_first_level_2__13__q  & ((Xd_0__inst_inst_first_level_0__13__q ) # 
// (Xd_0__inst_inst_first_level_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__13__q ),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_50 ),
	.sharein(Xd_0__inst_inst_inst_rtl_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_53_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_54 ),
	.shareout(Xd_0__inst_inst_inst_rtl_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_57 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_57_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__14__q  $ (!Xd_0__inst_inst_first_level_1__14__q  $ (Xd_0__inst_inst_first_level_0__14__q )) ) + ( Xd_0__inst_inst_inst_rtl_55  ) + ( Xd_0__inst_inst_inst_rtl_54  ))
// Xd_0__inst_inst_inst_rtl_58  = CARRY(( !Xd_0__inst_inst_first_level_2__14__q  $ (!Xd_0__inst_inst_first_level_1__14__q  $ (Xd_0__inst_inst_first_level_0__14__q )) ) + ( Xd_0__inst_inst_inst_rtl_55  ) + ( Xd_0__inst_inst_inst_rtl_54  ))
// Xd_0__inst_inst_inst_rtl_59  = SHARE((!Xd_0__inst_inst_first_level_2__14__q  & (Xd_0__inst_inst_first_level_1__14__q  & Xd_0__inst_inst_first_level_0__14__q )) # (Xd_0__inst_inst_first_level_2__14__q  & ((Xd_0__inst_inst_first_level_0__14__q ) # 
// (Xd_0__inst_inst_first_level_1__14__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__14__q ),
	.datac(!Xd_0__inst_inst_first_level_1__14__q ),
	.datad(!Xd_0__inst_inst_first_level_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_54 ),
	.sharein(Xd_0__inst_inst_inst_rtl_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_57_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_58 ),
	.shareout(Xd_0__inst_inst_inst_rtl_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_61 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_61_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_rtl_59  ) + ( Xd_0__inst_inst_inst_rtl_58  ))
// Xd_0__inst_inst_inst_rtl_62  = CARRY(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_rtl_59  ) + ( Xd_0__inst_inst_inst_rtl_58  ))
// Xd_0__inst_inst_inst_rtl_63  = SHARE((!Xd_0__inst_inst_first_level_2__15__q  & (Xd_0__inst_inst_first_level_1__15__q  & Xd_0__inst_inst_first_level_0__15__q )) # (Xd_0__inst_inst_first_level_2__15__q  & ((Xd_0__inst_inst_first_level_0__15__q ) # 
// (Xd_0__inst_inst_first_level_1__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__15__q ),
	.datac(!Xd_0__inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_58 ),
	.sharein(Xd_0__inst_inst_inst_rtl_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_61_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_62 ),
	.shareout(Xd_0__inst_inst_inst_rtl_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_65 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_65_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__16__q  $ (!Xd_0__inst_inst_first_level_1__16__q  $ (Xd_0__inst_inst_first_level_0__16__q )) ) + ( Xd_0__inst_inst_inst_rtl_63  ) + ( Xd_0__inst_inst_inst_rtl_62  ))
// Xd_0__inst_inst_inst_rtl_66  = CARRY(( !Xd_0__inst_inst_first_level_2__16__q  $ (!Xd_0__inst_inst_first_level_1__16__q  $ (Xd_0__inst_inst_first_level_0__16__q )) ) + ( Xd_0__inst_inst_inst_rtl_63  ) + ( Xd_0__inst_inst_inst_rtl_62  ))
// Xd_0__inst_inst_inst_rtl_67  = SHARE((!Xd_0__inst_inst_first_level_2__16__q  & (Xd_0__inst_inst_first_level_1__16__q  & Xd_0__inst_inst_first_level_0__16__q )) # (Xd_0__inst_inst_first_level_2__16__q  & ((Xd_0__inst_inst_first_level_0__16__q ) # 
// (Xd_0__inst_inst_first_level_1__16__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__16__q ),
	.datac(!Xd_0__inst_inst_first_level_1__16__q ),
	.datad(!Xd_0__inst_inst_first_level_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_62 ),
	.sharein(Xd_0__inst_inst_inst_rtl_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_65_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_66 ),
	.shareout(Xd_0__inst_inst_inst_rtl_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_69 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_69_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__17__q  $ (!Xd_0__inst_inst_first_level_1__17__q  $ (Xd_0__inst_inst_first_level_0__17__q )) ) + ( Xd_0__inst_inst_inst_rtl_67  ) + ( Xd_0__inst_inst_inst_rtl_66  ))
// Xd_0__inst_inst_inst_rtl_70  = CARRY(( !Xd_0__inst_inst_first_level_2__17__q  $ (!Xd_0__inst_inst_first_level_1__17__q  $ (Xd_0__inst_inst_first_level_0__17__q )) ) + ( Xd_0__inst_inst_inst_rtl_67  ) + ( Xd_0__inst_inst_inst_rtl_66  ))
// Xd_0__inst_inst_inst_rtl_71  = SHARE((!Xd_0__inst_inst_first_level_2__17__q  & (Xd_0__inst_inst_first_level_1__17__q  & Xd_0__inst_inst_first_level_0__17__q )) # (Xd_0__inst_inst_first_level_2__17__q  & ((Xd_0__inst_inst_first_level_0__17__q ) # 
// (Xd_0__inst_inst_first_level_1__17__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__17__q ),
	.datac(!Xd_0__inst_inst_first_level_1__17__q ),
	.datad(!Xd_0__inst_inst_first_level_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_66 ),
	.sharein(Xd_0__inst_inst_inst_rtl_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_69_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_70 ),
	.shareout(Xd_0__inst_inst_inst_rtl_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_73 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_73_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__18__q  $ (!Xd_0__inst_inst_first_level_1__18__q  $ (Xd_0__inst_inst_first_level_0__18__q )) ) + ( Xd_0__inst_inst_inst_rtl_71  ) + ( Xd_0__inst_inst_inst_rtl_70  ))
// Xd_0__inst_inst_inst_rtl_74  = CARRY(( !Xd_0__inst_inst_first_level_2__18__q  $ (!Xd_0__inst_inst_first_level_1__18__q  $ (Xd_0__inst_inst_first_level_0__18__q )) ) + ( Xd_0__inst_inst_inst_rtl_71  ) + ( Xd_0__inst_inst_inst_rtl_70  ))
// Xd_0__inst_inst_inst_rtl_75  = SHARE((!Xd_0__inst_inst_first_level_2__18__q  & (Xd_0__inst_inst_first_level_1__18__q  & Xd_0__inst_inst_first_level_0__18__q )) # (Xd_0__inst_inst_first_level_2__18__q  & ((Xd_0__inst_inst_first_level_0__18__q ) # 
// (Xd_0__inst_inst_first_level_1__18__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__18__q ),
	.datac(!Xd_0__inst_inst_first_level_1__18__q ),
	.datad(!Xd_0__inst_inst_first_level_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_70 ),
	.sharein(Xd_0__inst_inst_inst_rtl_71 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_73_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_74 ),
	.shareout(Xd_0__inst_inst_inst_rtl_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_77 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_77_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__19__q  $ (!Xd_0__inst_inst_first_level_1__19__q  $ (Xd_0__inst_inst_first_level_0__19__q )) ) + ( Xd_0__inst_inst_inst_rtl_75  ) + ( Xd_0__inst_inst_inst_rtl_74  ))
// Xd_0__inst_inst_inst_rtl_78  = CARRY(( !Xd_0__inst_inst_first_level_2__19__q  $ (!Xd_0__inst_inst_first_level_1__19__q  $ (Xd_0__inst_inst_first_level_0__19__q )) ) + ( Xd_0__inst_inst_inst_rtl_75  ) + ( Xd_0__inst_inst_inst_rtl_74  ))
// Xd_0__inst_inst_inst_rtl_79  = SHARE((!Xd_0__inst_inst_first_level_2__19__q  & (Xd_0__inst_inst_first_level_1__19__q  & Xd_0__inst_inst_first_level_0__19__q )) # (Xd_0__inst_inst_first_level_2__19__q  & ((Xd_0__inst_inst_first_level_0__19__q ) # 
// (Xd_0__inst_inst_first_level_1__19__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__19__q ),
	.datac(!Xd_0__inst_inst_first_level_1__19__q ),
	.datad(!Xd_0__inst_inst_first_level_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_74 ),
	.sharein(Xd_0__inst_inst_inst_rtl_75 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_77_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_78 ),
	.shareout(Xd_0__inst_inst_inst_rtl_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_81 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_81_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__20__q  $ (!Xd_0__inst_inst_first_level_1__20__q  $ (Xd_0__inst_inst_first_level_0__20__q )) ) + ( Xd_0__inst_inst_inst_rtl_79  ) + ( Xd_0__inst_inst_inst_rtl_78  ))
// Xd_0__inst_inst_inst_rtl_82  = CARRY(( !Xd_0__inst_inst_first_level_2__20__q  $ (!Xd_0__inst_inst_first_level_1__20__q  $ (Xd_0__inst_inst_first_level_0__20__q )) ) + ( Xd_0__inst_inst_inst_rtl_79  ) + ( Xd_0__inst_inst_inst_rtl_78  ))
// Xd_0__inst_inst_inst_rtl_83  = SHARE((!Xd_0__inst_inst_first_level_2__20__q  & (Xd_0__inst_inst_first_level_1__20__q  & Xd_0__inst_inst_first_level_0__20__q )) # (Xd_0__inst_inst_first_level_2__20__q  & ((Xd_0__inst_inst_first_level_0__20__q ) # 
// (Xd_0__inst_inst_first_level_1__20__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__20__q ),
	.datac(!Xd_0__inst_inst_first_level_1__20__q ),
	.datad(!Xd_0__inst_inst_first_level_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_78 ),
	.sharein(Xd_0__inst_inst_inst_rtl_79 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_81_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_82 ),
	.shareout(Xd_0__inst_inst_inst_rtl_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_85 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_85_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__21__q  $ (!Xd_0__inst_inst_first_level_1__21__q  $ (Xd_0__inst_inst_first_level_0__21__q )) ) + ( Xd_0__inst_inst_inst_rtl_83  ) + ( Xd_0__inst_inst_inst_rtl_82  ))
// Xd_0__inst_inst_inst_rtl_86  = CARRY(( !Xd_0__inst_inst_first_level_2__21__q  $ (!Xd_0__inst_inst_first_level_1__21__q  $ (Xd_0__inst_inst_first_level_0__21__q )) ) + ( Xd_0__inst_inst_inst_rtl_83  ) + ( Xd_0__inst_inst_inst_rtl_82  ))
// Xd_0__inst_inst_inst_rtl_87  = SHARE((!Xd_0__inst_inst_first_level_2__21__q  & (Xd_0__inst_inst_first_level_1__21__q  & Xd_0__inst_inst_first_level_0__21__q )) # (Xd_0__inst_inst_first_level_2__21__q  & ((Xd_0__inst_inst_first_level_0__21__q ) # 
// (Xd_0__inst_inst_first_level_1__21__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__21__q ),
	.datac(!Xd_0__inst_inst_first_level_1__21__q ),
	.datad(!Xd_0__inst_inst_first_level_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_82 ),
	.sharein(Xd_0__inst_inst_inst_rtl_83 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_85_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_86 ),
	.shareout(Xd_0__inst_inst_inst_rtl_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_89 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_89_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__22__q  $ (!Xd_0__inst_inst_first_level_1__22__q  $ (Xd_0__inst_inst_first_level_0__22__q )) ) + ( Xd_0__inst_inst_inst_rtl_87  ) + ( Xd_0__inst_inst_inst_rtl_86  ))
// Xd_0__inst_inst_inst_rtl_90  = CARRY(( !Xd_0__inst_inst_first_level_2__22__q  $ (!Xd_0__inst_inst_first_level_1__22__q  $ (Xd_0__inst_inst_first_level_0__22__q )) ) + ( Xd_0__inst_inst_inst_rtl_87  ) + ( Xd_0__inst_inst_inst_rtl_86  ))
// Xd_0__inst_inst_inst_rtl_91  = SHARE((!Xd_0__inst_inst_first_level_2__22__q  & (Xd_0__inst_inst_first_level_1__22__q  & Xd_0__inst_inst_first_level_0__22__q )) # (Xd_0__inst_inst_first_level_2__22__q  & ((Xd_0__inst_inst_first_level_0__22__q ) # 
// (Xd_0__inst_inst_first_level_1__22__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__22__q ),
	.datac(!Xd_0__inst_inst_first_level_1__22__q ),
	.datad(!Xd_0__inst_inst_first_level_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_86 ),
	.sharein(Xd_0__inst_inst_inst_rtl_87 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_89_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_90 ),
	.shareout(Xd_0__inst_inst_inst_rtl_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_93 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_93_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__23__q  $ (!Xd_0__inst_inst_first_level_1__23__q  $ (Xd_0__inst_inst_first_level_0__23__q )) ) + ( Xd_0__inst_inst_inst_rtl_91  ) + ( Xd_0__inst_inst_inst_rtl_90  ))
// Xd_0__inst_inst_inst_rtl_94  = CARRY(( !Xd_0__inst_inst_first_level_2__23__q  $ (!Xd_0__inst_inst_first_level_1__23__q  $ (Xd_0__inst_inst_first_level_0__23__q )) ) + ( Xd_0__inst_inst_inst_rtl_91  ) + ( Xd_0__inst_inst_inst_rtl_90  ))
// Xd_0__inst_inst_inst_rtl_95  = SHARE((!Xd_0__inst_inst_first_level_2__23__q  & (Xd_0__inst_inst_first_level_1__23__q  & Xd_0__inst_inst_first_level_0__23__q )) # (Xd_0__inst_inst_first_level_2__23__q  & ((Xd_0__inst_inst_first_level_0__23__q ) # 
// (Xd_0__inst_inst_first_level_1__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__23__q ),
	.datac(!Xd_0__inst_inst_first_level_1__23__q ),
	.datad(!Xd_0__inst_inst_first_level_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_90 ),
	.sharein(Xd_0__inst_inst_inst_rtl_91 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_93_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_94 ),
	.shareout(Xd_0__inst_inst_inst_rtl_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_97 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_97_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__25__q  $ (!Xd_0__inst_inst_first_level_1__24__q  $ (Xd_0__inst_inst_first_level_0__24__q )) ) + ( Xd_0__inst_inst_inst_rtl_95  ) + ( Xd_0__inst_inst_inst_rtl_94  ))
// Xd_0__inst_inst_inst_rtl_98  = CARRY(( !Xd_0__inst_inst_first_level_2__25__q  $ (!Xd_0__inst_inst_first_level_1__24__q  $ (Xd_0__inst_inst_first_level_0__24__q )) ) + ( Xd_0__inst_inst_inst_rtl_95  ) + ( Xd_0__inst_inst_inst_rtl_94  ))
// Xd_0__inst_inst_inst_rtl_99  = SHARE((!Xd_0__inst_inst_first_level_2__25__q  & (Xd_0__inst_inst_first_level_1__24__q  & Xd_0__inst_inst_first_level_0__24__q )) # (Xd_0__inst_inst_first_level_2__25__q  & ((Xd_0__inst_inst_first_level_0__24__q ) # 
// (Xd_0__inst_inst_first_level_1__24__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__25__q ),
	.datac(!Xd_0__inst_inst_first_level_1__24__q ),
	.datad(!Xd_0__inst_inst_first_level_0__24__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_94 ),
	.sharein(Xd_0__inst_inst_inst_rtl_95 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_97_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_98 ),
	.shareout(Xd_0__inst_inst_inst_rtl_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_101 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_101_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__25__q  $ (!Xd_0__inst_inst_first_level_1__25__q  $ (Xd_0__inst_inst_first_level_0__25__q )) ) + ( Xd_0__inst_inst_inst_rtl_99  ) + ( Xd_0__inst_inst_inst_rtl_98  ))
// Xd_0__inst_inst_inst_rtl_102  = CARRY(( !Xd_0__inst_inst_first_level_2__25__q  $ (!Xd_0__inst_inst_first_level_1__25__q  $ (Xd_0__inst_inst_first_level_0__25__q )) ) + ( Xd_0__inst_inst_inst_rtl_99  ) + ( Xd_0__inst_inst_inst_rtl_98  ))
// Xd_0__inst_inst_inst_rtl_103  = SHARE((!Xd_0__inst_inst_first_level_2__25__q  & (Xd_0__inst_inst_first_level_1__25__q  & Xd_0__inst_inst_first_level_0__25__q )) # (Xd_0__inst_inst_first_level_2__25__q  & ((Xd_0__inst_inst_first_level_0__25__q ) # 
// (Xd_0__inst_inst_first_level_1__25__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__25__q ),
	.datac(!Xd_0__inst_inst_first_level_1__25__q ),
	.datad(!Xd_0__inst_inst_first_level_0__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_98 ),
	.sharein(Xd_0__inst_inst_inst_rtl_99 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_101_sumout ),
	.cout(Xd_0__inst_inst_inst_rtl_102 ),
	.shareout(Xd_0__inst_inst_inst_rtl_103 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_rtl_105 (
// Equation(s):
// Xd_0__inst_inst_inst_rtl_105_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__25__q  $ (!Xd_0__inst_inst_first_level_1__25__q  $ (Xd_0__inst_inst_first_level_0__25__q )) ) + ( Xd_0__inst_inst_inst_rtl_103  ) + ( Xd_0__inst_inst_inst_rtl_102  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__25__q ),
	.datac(!Xd_0__inst_inst_first_level_1__25__q ),
	.datad(!Xd_0__inst_inst_first_level_0__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_rtl_102 ),
	.sharein(Xd_0__inst_inst_inst_rtl_103 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_rtl_105_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_172 (
// Equation(s):
// Xd_0__inst_mult_4_173  = SUM(( GND ) + ( Xd_0__inst_mult_4_179  ) + ( Xd_0__inst_mult_4_178  ))
// Xd_0__inst_mult_4_174  = CARRY(( GND ) + ( Xd_0__inst_mult_4_179  ) + ( Xd_0__inst_mult_4_178  ))
// Xd_0__inst_mult_4_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_178 ),
	.sharein(Xd_0__inst_mult_4_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_173 ),
	.cout(Xd_0__inst_mult_4_174 ),
	.shareout(Xd_0__inst_mult_4_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_1 (
// Equation(s):
// Xd_0__inst_inst_add_4_1_sumout  = SUM(( !Xd_0__inst_r_sum1_6__0__q  $ (!Xd_0__inst_r_sum1_7__0__q ) ) + ( Xd_0__inst_mult_14_175  ) + ( Xd_0__inst_mult_14_174  ))
// Xd_0__inst_inst_add_4_2  = CARRY(( !Xd_0__inst_r_sum1_6__0__q  $ (!Xd_0__inst_r_sum1_7__0__q ) ) + ( Xd_0__inst_mult_14_175  ) + ( Xd_0__inst_mult_14_174  ))
// Xd_0__inst_inst_add_4_3  = SHARE((Xd_0__inst_r_sum1_6__0__q  & Xd_0__inst_r_sum1_7__0__q ))

	.dataa(!Xd_0__inst_r_sum1_6__0__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_174 ),
	.sharein(Xd_0__inst_mult_14_175 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_1_sumout ),
	.cout(Xd_0__inst_inst_add_4_2 ),
	.shareout(Xd_0__inst_inst_add_4_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_1 (
// Equation(s):
// Xd_0__inst_inst_add_2_1_sumout  = SUM(( !Xd_0__inst_r_sum1_5__0__q  $ (!Xd_0__inst_r_sum1_4__0__q  $ (Xd_0__inst_r_sum1_3__0__q )) ) + ( Xd_0__inst_mult_15_175  ) + ( Xd_0__inst_mult_15_174  ))
// Xd_0__inst_inst_add_2_2  = CARRY(( !Xd_0__inst_r_sum1_5__0__q  $ (!Xd_0__inst_r_sum1_4__0__q  $ (Xd_0__inst_r_sum1_3__0__q )) ) + ( Xd_0__inst_mult_15_175  ) + ( Xd_0__inst_mult_15_174  ))
// Xd_0__inst_inst_add_2_3  = SHARE((!Xd_0__inst_r_sum1_5__0__q  & (Xd_0__inst_r_sum1_4__0__q  & Xd_0__inst_r_sum1_3__0__q )) # (Xd_0__inst_r_sum1_5__0__q  & ((Xd_0__inst_r_sum1_3__0__q ) # (Xd_0__inst_r_sum1_4__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__0__q ),
	.datac(!Xd_0__inst_r_sum1_4__0__q ),
	.datad(!Xd_0__inst_r_sum1_3__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_174 ),
	.sharein(Xd_0__inst_mult_15_175 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_1_sumout ),
	.cout(Xd_0__inst_inst_add_2_2 ),
	.shareout(Xd_0__inst_inst_add_2_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_mult_12_171  ) + ( Xd_0__inst_mult_12_170  ))
// Xd_0__inst_inst_add_0_2  = CARRY(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_mult_12_171  ) + ( Xd_0__inst_mult_12_170  ))
// Xd_0__inst_inst_add_0_3  = SHARE((!Xd_0__inst_r_sum1_2__0__q  & (Xd_0__inst_r_sum1_1__0__q  & Xd_0__inst_r_sum1_0__0__q )) # (Xd_0__inst_r_sum1_2__0__q  & ((Xd_0__inst_r_sum1_0__0__q ) # (Xd_0__inst_r_sum1_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__0__q ),
	.datac(!Xd_0__inst_r_sum1_1__0__q ),
	.datad(!Xd_0__inst_r_sum1_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_170 ),
	.sharein(Xd_0__inst_mult_12_171 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4 (
// Equation(s):
// Xd_0__inst_mult_4_177  = SUM(( (din_a[56] & din_b[58]) ) + ( Xd_0__inst_mult_4_182  ) + ( Xd_0__inst_mult_4_181  ))
// Xd_0__inst_mult_4_178  = CARRY(( (din_a[56] & din_b[58]) ) + ( Xd_0__inst_mult_4_182  ) + ( Xd_0__inst_mult_4_181  ))
// Xd_0__inst_mult_4_179  = SHARE(GND)

	.dataa(!din_a[56]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_181 ),
	.sharein(Xd_0__inst_mult_4_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_177 ),
	.cout(Xd_0__inst_mult_4_178 ),
	.shareout(Xd_0__inst_mult_4_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_5 (
// Equation(s):
// Xd_0__inst_inst_add_4_5_sumout  = SUM(( !Xd_0__inst_r_sum1_6__1__q  $ (!Xd_0__inst_r_sum1_7__1__q ) ) + ( Xd_0__inst_inst_add_4_3  ) + ( Xd_0__inst_inst_add_4_2  ))
// Xd_0__inst_inst_add_4_6  = CARRY(( !Xd_0__inst_r_sum1_6__1__q  $ (!Xd_0__inst_r_sum1_7__1__q ) ) + ( Xd_0__inst_inst_add_4_3  ) + ( Xd_0__inst_inst_add_4_2  ))
// Xd_0__inst_inst_add_4_7  = SHARE((Xd_0__inst_r_sum1_6__1__q  & Xd_0__inst_r_sum1_7__1__q ))

	.dataa(!Xd_0__inst_r_sum1_6__1__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_2 ),
	.sharein(Xd_0__inst_inst_add_4_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_5_sumout ),
	.cout(Xd_0__inst_inst_add_4_6 ),
	.shareout(Xd_0__inst_inst_add_4_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_5 (
// Equation(s):
// Xd_0__inst_inst_add_2_5_sumout  = SUM(( !Xd_0__inst_r_sum1_5__1__q  $ (!Xd_0__inst_r_sum1_4__1__q  $ (Xd_0__inst_r_sum1_3__1__q )) ) + ( Xd_0__inst_inst_add_2_3  ) + ( Xd_0__inst_inst_add_2_2  ))
// Xd_0__inst_inst_add_2_6  = CARRY(( !Xd_0__inst_r_sum1_5__1__q  $ (!Xd_0__inst_r_sum1_4__1__q  $ (Xd_0__inst_r_sum1_3__1__q )) ) + ( Xd_0__inst_inst_add_2_3  ) + ( Xd_0__inst_inst_add_2_2  ))
// Xd_0__inst_inst_add_2_7  = SHARE((!Xd_0__inst_r_sum1_5__1__q  & (Xd_0__inst_r_sum1_4__1__q  & Xd_0__inst_r_sum1_3__1__q )) # (Xd_0__inst_r_sum1_5__1__q  & ((Xd_0__inst_r_sum1_3__1__q ) # (Xd_0__inst_r_sum1_4__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__1__q ),
	.datac(!Xd_0__inst_r_sum1_4__1__q ),
	.datad(!Xd_0__inst_r_sum1_3__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_2 ),
	.sharein(Xd_0__inst_inst_add_2_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_5_sumout ),
	.cout(Xd_0__inst_inst_add_2_6 ),
	.shareout(Xd_0__inst_inst_add_2_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_6  = CARRY(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_7  = SHARE((!Xd_0__inst_r_sum1_2__1__q  & (Xd_0__inst_r_sum1_1__1__q  & Xd_0__inst_r_sum1_0__1__q )) # (Xd_0__inst_r_sum1_2__1__q  & ((Xd_0__inst_r_sum1_0__1__q ) # (Xd_0__inst_r_sum1_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__1__q ),
	.datac(!Xd_0__inst_r_sum1_1__1__q ),
	.datad(!Xd_0__inst_r_sum1_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_9 (
// Equation(s):
// Xd_0__inst_inst_add_4_9_sumout  = SUM(( !Xd_0__inst_r_sum1_6__2__q  $ (!Xd_0__inst_r_sum1_7__2__q ) ) + ( Xd_0__inst_inst_add_4_7  ) + ( Xd_0__inst_inst_add_4_6  ))
// Xd_0__inst_inst_add_4_10  = CARRY(( !Xd_0__inst_r_sum1_6__2__q  $ (!Xd_0__inst_r_sum1_7__2__q ) ) + ( Xd_0__inst_inst_add_4_7  ) + ( Xd_0__inst_inst_add_4_6  ))
// Xd_0__inst_inst_add_4_11  = SHARE((Xd_0__inst_r_sum1_6__2__q  & Xd_0__inst_r_sum1_7__2__q ))

	.dataa(!Xd_0__inst_r_sum1_6__2__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_6 ),
	.sharein(Xd_0__inst_inst_add_4_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_9_sumout ),
	.cout(Xd_0__inst_inst_add_4_10 ),
	.shareout(Xd_0__inst_inst_add_4_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_9 (
// Equation(s):
// Xd_0__inst_inst_add_2_9_sumout  = SUM(( !Xd_0__inst_r_sum1_5__2__q  $ (!Xd_0__inst_r_sum1_4__2__q  $ (Xd_0__inst_r_sum1_3__2__q )) ) + ( Xd_0__inst_inst_add_2_7  ) + ( Xd_0__inst_inst_add_2_6  ))
// Xd_0__inst_inst_add_2_10  = CARRY(( !Xd_0__inst_r_sum1_5__2__q  $ (!Xd_0__inst_r_sum1_4__2__q  $ (Xd_0__inst_r_sum1_3__2__q )) ) + ( Xd_0__inst_inst_add_2_7  ) + ( Xd_0__inst_inst_add_2_6  ))
// Xd_0__inst_inst_add_2_11  = SHARE((!Xd_0__inst_r_sum1_5__2__q  & (Xd_0__inst_r_sum1_4__2__q  & Xd_0__inst_r_sum1_3__2__q )) # (Xd_0__inst_r_sum1_5__2__q  & ((Xd_0__inst_r_sum1_3__2__q ) # (Xd_0__inst_r_sum1_4__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__2__q ),
	.datac(!Xd_0__inst_r_sum1_4__2__q ),
	.datad(!Xd_0__inst_r_sum1_3__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_6 ),
	.sharein(Xd_0__inst_inst_add_2_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_9_sumout ),
	.cout(Xd_0__inst_inst_add_2_10 ),
	.shareout(Xd_0__inst_inst_add_2_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_10  = CARRY(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_11  = SHARE((!Xd_0__inst_r_sum1_2__2__q  & (Xd_0__inst_r_sum1_1__2__q  & Xd_0__inst_r_sum1_0__2__q )) # (Xd_0__inst_r_sum1_2__2__q  & ((Xd_0__inst_r_sum1_0__2__q ) # (Xd_0__inst_r_sum1_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__2__q ),
	.datac(!Xd_0__inst_r_sum1_1__2__q ),
	.datad(!Xd_0__inst_r_sum1_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_13 (
// Equation(s):
// Xd_0__inst_inst_add_4_13_sumout  = SUM(( !Xd_0__inst_r_sum1_6__3__q  $ (!Xd_0__inst_r_sum1_7__3__q ) ) + ( Xd_0__inst_inst_add_4_11  ) + ( Xd_0__inst_inst_add_4_10  ))
// Xd_0__inst_inst_add_4_14  = CARRY(( !Xd_0__inst_r_sum1_6__3__q  $ (!Xd_0__inst_r_sum1_7__3__q ) ) + ( Xd_0__inst_inst_add_4_11  ) + ( Xd_0__inst_inst_add_4_10  ))
// Xd_0__inst_inst_add_4_15  = SHARE((Xd_0__inst_r_sum1_6__3__q  & Xd_0__inst_r_sum1_7__3__q ))

	.dataa(!Xd_0__inst_r_sum1_6__3__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_10 ),
	.sharein(Xd_0__inst_inst_add_4_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_13_sumout ),
	.cout(Xd_0__inst_inst_add_4_14 ),
	.shareout(Xd_0__inst_inst_add_4_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_13 (
// Equation(s):
// Xd_0__inst_inst_add_2_13_sumout  = SUM(( !Xd_0__inst_r_sum1_5__3__q  $ (!Xd_0__inst_r_sum1_4__3__q  $ (Xd_0__inst_r_sum1_3__3__q )) ) + ( Xd_0__inst_inst_add_2_11  ) + ( Xd_0__inst_inst_add_2_10  ))
// Xd_0__inst_inst_add_2_14  = CARRY(( !Xd_0__inst_r_sum1_5__3__q  $ (!Xd_0__inst_r_sum1_4__3__q  $ (Xd_0__inst_r_sum1_3__3__q )) ) + ( Xd_0__inst_inst_add_2_11  ) + ( Xd_0__inst_inst_add_2_10  ))
// Xd_0__inst_inst_add_2_15  = SHARE((!Xd_0__inst_r_sum1_5__3__q  & (Xd_0__inst_r_sum1_4__3__q  & Xd_0__inst_r_sum1_3__3__q )) # (Xd_0__inst_r_sum1_5__3__q  & ((Xd_0__inst_r_sum1_3__3__q ) # (Xd_0__inst_r_sum1_4__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__3__q ),
	.datac(!Xd_0__inst_r_sum1_4__3__q ),
	.datad(!Xd_0__inst_r_sum1_3__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_10 ),
	.sharein(Xd_0__inst_inst_add_2_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_13_sumout ),
	.cout(Xd_0__inst_inst_add_2_14 ),
	.shareout(Xd_0__inst_inst_add_2_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_14  = CARRY(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_15  = SHARE((!Xd_0__inst_r_sum1_2__3__q  & (Xd_0__inst_r_sum1_1__3__q  & Xd_0__inst_r_sum1_0__3__q )) # (Xd_0__inst_r_sum1_2__3__q  & ((Xd_0__inst_r_sum1_0__3__q ) # (Xd_0__inst_r_sum1_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__3__q ),
	.datac(!Xd_0__inst_r_sum1_1__3__q ),
	.datad(!Xd_0__inst_r_sum1_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_17 (
// Equation(s):
// Xd_0__inst_inst_add_4_17_sumout  = SUM(( !Xd_0__inst_r_sum1_6__4__q  $ (!Xd_0__inst_r_sum1_7__4__q ) ) + ( Xd_0__inst_inst_add_4_15  ) + ( Xd_0__inst_inst_add_4_14  ))
// Xd_0__inst_inst_add_4_18  = CARRY(( !Xd_0__inst_r_sum1_6__4__q  $ (!Xd_0__inst_r_sum1_7__4__q ) ) + ( Xd_0__inst_inst_add_4_15  ) + ( Xd_0__inst_inst_add_4_14  ))
// Xd_0__inst_inst_add_4_19  = SHARE((Xd_0__inst_r_sum1_6__4__q  & Xd_0__inst_r_sum1_7__4__q ))

	.dataa(!Xd_0__inst_r_sum1_6__4__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_14 ),
	.sharein(Xd_0__inst_inst_add_4_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_17_sumout ),
	.cout(Xd_0__inst_inst_add_4_18 ),
	.shareout(Xd_0__inst_inst_add_4_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_17 (
// Equation(s):
// Xd_0__inst_inst_add_2_17_sumout  = SUM(( !Xd_0__inst_r_sum1_5__4__q  $ (!Xd_0__inst_r_sum1_4__4__q  $ (Xd_0__inst_r_sum1_3__4__q )) ) + ( Xd_0__inst_inst_add_2_15  ) + ( Xd_0__inst_inst_add_2_14  ))
// Xd_0__inst_inst_add_2_18  = CARRY(( !Xd_0__inst_r_sum1_5__4__q  $ (!Xd_0__inst_r_sum1_4__4__q  $ (Xd_0__inst_r_sum1_3__4__q )) ) + ( Xd_0__inst_inst_add_2_15  ) + ( Xd_0__inst_inst_add_2_14  ))
// Xd_0__inst_inst_add_2_19  = SHARE((!Xd_0__inst_r_sum1_5__4__q  & (Xd_0__inst_r_sum1_4__4__q  & Xd_0__inst_r_sum1_3__4__q )) # (Xd_0__inst_r_sum1_5__4__q  & ((Xd_0__inst_r_sum1_3__4__q ) # (Xd_0__inst_r_sum1_4__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__4__q ),
	.datac(!Xd_0__inst_r_sum1_4__4__q ),
	.datad(!Xd_0__inst_r_sum1_3__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_14 ),
	.sharein(Xd_0__inst_inst_add_2_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_17_sumout ),
	.cout(Xd_0__inst_inst_add_2_18 ),
	.shareout(Xd_0__inst_inst_add_2_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_18  = CARRY(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_19  = SHARE((!Xd_0__inst_r_sum1_2__4__q  & (Xd_0__inst_r_sum1_1__4__q  & Xd_0__inst_r_sum1_0__4__q )) # (Xd_0__inst_r_sum1_2__4__q  & ((Xd_0__inst_r_sum1_0__4__q ) # (Xd_0__inst_r_sum1_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__4__q ),
	.datac(!Xd_0__inst_r_sum1_1__4__q ),
	.datad(!Xd_0__inst_r_sum1_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_21 (
// Equation(s):
// Xd_0__inst_inst_add_4_21_sumout  = SUM(( !Xd_0__inst_r_sum1_6__5__q  $ (!Xd_0__inst_r_sum1_7__5__q ) ) + ( Xd_0__inst_inst_add_4_19  ) + ( Xd_0__inst_inst_add_4_18  ))
// Xd_0__inst_inst_add_4_22  = CARRY(( !Xd_0__inst_r_sum1_6__5__q  $ (!Xd_0__inst_r_sum1_7__5__q ) ) + ( Xd_0__inst_inst_add_4_19  ) + ( Xd_0__inst_inst_add_4_18  ))
// Xd_0__inst_inst_add_4_23  = SHARE((Xd_0__inst_r_sum1_6__5__q  & Xd_0__inst_r_sum1_7__5__q ))

	.dataa(!Xd_0__inst_r_sum1_6__5__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_18 ),
	.sharein(Xd_0__inst_inst_add_4_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_21_sumout ),
	.cout(Xd_0__inst_inst_add_4_22 ),
	.shareout(Xd_0__inst_inst_add_4_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_21 (
// Equation(s):
// Xd_0__inst_inst_add_2_21_sumout  = SUM(( !Xd_0__inst_r_sum1_5__5__q  $ (!Xd_0__inst_r_sum1_4__5__q  $ (Xd_0__inst_r_sum1_3__5__q )) ) + ( Xd_0__inst_inst_add_2_19  ) + ( Xd_0__inst_inst_add_2_18  ))
// Xd_0__inst_inst_add_2_22  = CARRY(( !Xd_0__inst_r_sum1_5__5__q  $ (!Xd_0__inst_r_sum1_4__5__q  $ (Xd_0__inst_r_sum1_3__5__q )) ) + ( Xd_0__inst_inst_add_2_19  ) + ( Xd_0__inst_inst_add_2_18  ))
// Xd_0__inst_inst_add_2_23  = SHARE((!Xd_0__inst_r_sum1_5__5__q  & (Xd_0__inst_r_sum1_4__5__q  & Xd_0__inst_r_sum1_3__5__q )) # (Xd_0__inst_r_sum1_5__5__q  & ((Xd_0__inst_r_sum1_3__5__q ) # (Xd_0__inst_r_sum1_4__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__5__q ),
	.datac(!Xd_0__inst_r_sum1_4__5__q ),
	.datad(!Xd_0__inst_r_sum1_3__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_18 ),
	.sharein(Xd_0__inst_inst_add_2_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_21_sumout ),
	.cout(Xd_0__inst_inst_add_2_22 ),
	.shareout(Xd_0__inst_inst_add_2_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_22  = CARRY(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_23  = SHARE((!Xd_0__inst_r_sum1_2__5__q  & (Xd_0__inst_r_sum1_1__5__q  & Xd_0__inst_r_sum1_0__5__q )) # (Xd_0__inst_r_sum1_2__5__q  & ((Xd_0__inst_r_sum1_0__5__q ) # (Xd_0__inst_r_sum1_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__5__q ),
	.datac(!Xd_0__inst_r_sum1_1__5__q ),
	.datad(!Xd_0__inst_r_sum1_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_25 (
// Equation(s):
// Xd_0__inst_inst_add_4_25_sumout  = SUM(( !Xd_0__inst_r_sum1_6__6__q  $ (!Xd_0__inst_r_sum1_7__6__q ) ) + ( Xd_0__inst_inst_add_4_23  ) + ( Xd_0__inst_inst_add_4_22  ))
// Xd_0__inst_inst_add_4_26  = CARRY(( !Xd_0__inst_r_sum1_6__6__q  $ (!Xd_0__inst_r_sum1_7__6__q ) ) + ( Xd_0__inst_inst_add_4_23  ) + ( Xd_0__inst_inst_add_4_22  ))
// Xd_0__inst_inst_add_4_27  = SHARE((Xd_0__inst_r_sum1_6__6__q  & Xd_0__inst_r_sum1_7__6__q ))

	.dataa(!Xd_0__inst_r_sum1_6__6__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_22 ),
	.sharein(Xd_0__inst_inst_add_4_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_25_sumout ),
	.cout(Xd_0__inst_inst_add_4_26 ),
	.shareout(Xd_0__inst_inst_add_4_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_25 (
// Equation(s):
// Xd_0__inst_inst_add_2_25_sumout  = SUM(( !Xd_0__inst_r_sum1_5__6__q  $ (!Xd_0__inst_r_sum1_4__6__q  $ (Xd_0__inst_r_sum1_3__6__q )) ) + ( Xd_0__inst_inst_add_2_23  ) + ( Xd_0__inst_inst_add_2_22  ))
// Xd_0__inst_inst_add_2_26  = CARRY(( !Xd_0__inst_r_sum1_5__6__q  $ (!Xd_0__inst_r_sum1_4__6__q  $ (Xd_0__inst_r_sum1_3__6__q )) ) + ( Xd_0__inst_inst_add_2_23  ) + ( Xd_0__inst_inst_add_2_22  ))
// Xd_0__inst_inst_add_2_27  = SHARE((!Xd_0__inst_r_sum1_5__6__q  & (Xd_0__inst_r_sum1_4__6__q  & Xd_0__inst_r_sum1_3__6__q )) # (Xd_0__inst_r_sum1_5__6__q  & ((Xd_0__inst_r_sum1_3__6__q ) # (Xd_0__inst_r_sum1_4__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__6__q ),
	.datac(!Xd_0__inst_r_sum1_4__6__q ),
	.datad(!Xd_0__inst_r_sum1_3__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_22 ),
	.sharein(Xd_0__inst_inst_add_2_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_25_sumout ),
	.cout(Xd_0__inst_inst_add_2_26 ),
	.shareout(Xd_0__inst_inst_add_2_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_26  = CARRY(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_27  = SHARE((!Xd_0__inst_r_sum1_2__6__q  & (Xd_0__inst_r_sum1_1__6__q  & Xd_0__inst_r_sum1_0__6__q )) # (Xd_0__inst_r_sum1_2__6__q  & ((Xd_0__inst_r_sum1_0__6__q ) # (Xd_0__inst_r_sum1_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__6__q ),
	.datac(!Xd_0__inst_r_sum1_1__6__q ),
	.datad(!Xd_0__inst_r_sum1_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_29 (
// Equation(s):
// Xd_0__inst_inst_add_4_29_sumout  = SUM(( !Xd_0__inst_r_sum1_6__7__q  $ (!Xd_0__inst_r_sum1_7__7__q ) ) + ( Xd_0__inst_inst_add_4_27  ) + ( Xd_0__inst_inst_add_4_26  ))
// Xd_0__inst_inst_add_4_30  = CARRY(( !Xd_0__inst_r_sum1_6__7__q  $ (!Xd_0__inst_r_sum1_7__7__q ) ) + ( Xd_0__inst_inst_add_4_27  ) + ( Xd_0__inst_inst_add_4_26  ))
// Xd_0__inst_inst_add_4_31  = SHARE((Xd_0__inst_r_sum1_6__7__q  & Xd_0__inst_r_sum1_7__7__q ))

	.dataa(!Xd_0__inst_r_sum1_6__7__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_26 ),
	.sharein(Xd_0__inst_inst_add_4_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_29_sumout ),
	.cout(Xd_0__inst_inst_add_4_30 ),
	.shareout(Xd_0__inst_inst_add_4_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_29 (
// Equation(s):
// Xd_0__inst_inst_add_2_29_sumout  = SUM(( !Xd_0__inst_r_sum1_5__7__q  $ (!Xd_0__inst_r_sum1_4__7__q  $ (Xd_0__inst_r_sum1_3__7__q )) ) + ( Xd_0__inst_inst_add_2_27  ) + ( Xd_0__inst_inst_add_2_26  ))
// Xd_0__inst_inst_add_2_30  = CARRY(( !Xd_0__inst_r_sum1_5__7__q  $ (!Xd_0__inst_r_sum1_4__7__q  $ (Xd_0__inst_r_sum1_3__7__q )) ) + ( Xd_0__inst_inst_add_2_27  ) + ( Xd_0__inst_inst_add_2_26  ))
// Xd_0__inst_inst_add_2_31  = SHARE((!Xd_0__inst_r_sum1_5__7__q  & (Xd_0__inst_r_sum1_4__7__q  & Xd_0__inst_r_sum1_3__7__q )) # (Xd_0__inst_r_sum1_5__7__q  & ((Xd_0__inst_r_sum1_3__7__q ) # (Xd_0__inst_r_sum1_4__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__7__q ),
	.datac(!Xd_0__inst_r_sum1_4__7__q ),
	.datad(!Xd_0__inst_r_sum1_3__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_26 ),
	.sharein(Xd_0__inst_inst_add_2_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_29_sumout ),
	.cout(Xd_0__inst_inst_add_2_30 ),
	.shareout(Xd_0__inst_inst_add_2_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_30  = CARRY(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_31  = SHARE((!Xd_0__inst_r_sum1_2__7__q  & (Xd_0__inst_r_sum1_1__7__q  & Xd_0__inst_r_sum1_0__7__q )) # (Xd_0__inst_r_sum1_2__7__q  & ((Xd_0__inst_r_sum1_0__7__q ) # (Xd_0__inst_r_sum1_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__7__q ),
	.datac(!Xd_0__inst_r_sum1_1__7__q ),
	.datad(!Xd_0__inst_r_sum1_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_33 (
// Equation(s):
// Xd_0__inst_inst_add_4_33_sumout  = SUM(( !Xd_0__inst_r_sum1_6__8__q  $ (!Xd_0__inst_r_sum1_7__8__q ) ) + ( Xd_0__inst_inst_add_4_31  ) + ( Xd_0__inst_inst_add_4_30  ))
// Xd_0__inst_inst_add_4_34  = CARRY(( !Xd_0__inst_r_sum1_6__8__q  $ (!Xd_0__inst_r_sum1_7__8__q ) ) + ( Xd_0__inst_inst_add_4_31  ) + ( Xd_0__inst_inst_add_4_30  ))
// Xd_0__inst_inst_add_4_35  = SHARE((Xd_0__inst_r_sum1_6__8__q  & Xd_0__inst_r_sum1_7__8__q ))

	.dataa(!Xd_0__inst_r_sum1_6__8__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_30 ),
	.sharein(Xd_0__inst_inst_add_4_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_33_sumout ),
	.cout(Xd_0__inst_inst_add_4_34 ),
	.shareout(Xd_0__inst_inst_add_4_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_33 (
// Equation(s):
// Xd_0__inst_inst_add_2_33_sumout  = SUM(( !Xd_0__inst_r_sum1_5__8__q  $ (!Xd_0__inst_r_sum1_4__8__q  $ (Xd_0__inst_r_sum1_3__8__q )) ) + ( Xd_0__inst_inst_add_2_31  ) + ( Xd_0__inst_inst_add_2_30  ))
// Xd_0__inst_inst_add_2_34  = CARRY(( !Xd_0__inst_r_sum1_5__8__q  $ (!Xd_0__inst_r_sum1_4__8__q  $ (Xd_0__inst_r_sum1_3__8__q )) ) + ( Xd_0__inst_inst_add_2_31  ) + ( Xd_0__inst_inst_add_2_30  ))
// Xd_0__inst_inst_add_2_35  = SHARE((!Xd_0__inst_r_sum1_5__8__q  & (Xd_0__inst_r_sum1_4__8__q  & Xd_0__inst_r_sum1_3__8__q )) # (Xd_0__inst_r_sum1_5__8__q  & ((Xd_0__inst_r_sum1_3__8__q ) # (Xd_0__inst_r_sum1_4__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__8__q ),
	.datac(!Xd_0__inst_r_sum1_4__8__q ),
	.datad(!Xd_0__inst_r_sum1_3__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_30 ),
	.sharein(Xd_0__inst_inst_add_2_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_33_sumout ),
	.cout(Xd_0__inst_inst_add_2_34 ),
	.shareout(Xd_0__inst_inst_add_2_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_34  = CARRY(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_35  = SHARE((!Xd_0__inst_r_sum1_2__8__q  & (Xd_0__inst_r_sum1_1__8__q  & Xd_0__inst_r_sum1_0__8__q )) # (Xd_0__inst_r_sum1_2__8__q  & ((Xd_0__inst_r_sum1_0__8__q ) # (Xd_0__inst_r_sum1_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__8__q ),
	.datac(!Xd_0__inst_r_sum1_1__8__q ),
	.datad(!Xd_0__inst_r_sum1_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_37 (
// Equation(s):
// Xd_0__inst_inst_add_4_37_sumout  = SUM(( !Xd_0__inst_r_sum1_6__9__q  $ (!Xd_0__inst_r_sum1_7__9__q ) ) + ( Xd_0__inst_inst_add_4_35  ) + ( Xd_0__inst_inst_add_4_34  ))
// Xd_0__inst_inst_add_4_38  = CARRY(( !Xd_0__inst_r_sum1_6__9__q  $ (!Xd_0__inst_r_sum1_7__9__q ) ) + ( Xd_0__inst_inst_add_4_35  ) + ( Xd_0__inst_inst_add_4_34  ))
// Xd_0__inst_inst_add_4_39  = SHARE((Xd_0__inst_r_sum1_6__9__q  & Xd_0__inst_r_sum1_7__9__q ))

	.dataa(!Xd_0__inst_r_sum1_6__9__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_34 ),
	.sharein(Xd_0__inst_inst_add_4_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_37_sumout ),
	.cout(Xd_0__inst_inst_add_4_38 ),
	.shareout(Xd_0__inst_inst_add_4_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_37 (
// Equation(s):
// Xd_0__inst_inst_add_2_37_sumout  = SUM(( !Xd_0__inst_r_sum1_5__9__q  $ (!Xd_0__inst_r_sum1_4__9__q  $ (Xd_0__inst_r_sum1_3__9__q )) ) + ( Xd_0__inst_inst_add_2_35  ) + ( Xd_0__inst_inst_add_2_34  ))
// Xd_0__inst_inst_add_2_38  = CARRY(( !Xd_0__inst_r_sum1_5__9__q  $ (!Xd_0__inst_r_sum1_4__9__q  $ (Xd_0__inst_r_sum1_3__9__q )) ) + ( Xd_0__inst_inst_add_2_35  ) + ( Xd_0__inst_inst_add_2_34  ))
// Xd_0__inst_inst_add_2_39  = SHARE((!Xd_0__inst_r_sum1_5__9__q  & (Xd_0__inst_r_sum1_4__9__q  & Xd_0__inst_r_sum1_3__9__q )) # (Xd_0__inst_r_sum1_5__9__q  & ((Xd_0__inst_r_sum1_3__9__q ) # (Xd_0__inst_r_sum1_4__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__9__q ),
	.datac(!Xd_0__inst_r_sum1_4__9__q ),
	.datad(!Xd_0__inst_r_sum1_3__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_34 ),
	.sharein(Xd_0__inst_inst_add_2_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_37_sumout ),
	.cout(Xd_0__inst_inst_add_2_38 ),
	.shareout(Xd_0__inst_inst_add_2_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_38  = CARRY(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_39  = SHARE((!Xd_0__inst_r_sum1_2__9__q  & (Xd_0__inst_r_sum1_1__9__q  & Xd_0__inst_r_sum1_0__9__q )) # (Xd_0__inst_r_sum1_2__9__q  & ((Xd_0__inst_r_sum1_0__9__q ) # (Xd_0__inst_r_sum1_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__9__q ),
	.datac(!Xd_0__inst_r_sum1_1__9__q ),
	.datad(!Xd_0__inst_r_sum1_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_41 (
// Equation(s):
// Xd_0__inst_inst_add_4_41_sumout  = SUM(( !Xd_0__inst_r_sum1_6__10__q  $ (!Xd_0__inst_r_sum1_7__10__q ) ) + ( Xd_0__inst_inst_add_4_39  ) + ( Xd_0__inst_inst_add_4_38  ))
// Xd_0__inst_inst_add_4_42  = CARRY(( !Xd_0__inst_r_sum1_6__10__q  $ (!Xd_0__inst_r_sum1_7__10__q ) ) + ( Xd_0__inst_inst_add_4_39  ) + ( Xd_0__inst_inst_add_4_38  ))
// Xd_0__inst_inst_add_4_43  = SHARE((Xd_0__inst_r_sum1_6__10__q  & Xd_0__inst_r_sum1_7__10__q ))

	.dataa(!Xd_0__inst_r_sum1_6__10__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_38 ),
	.sharein(Xd_0__inst_inst_add_4_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_41_sumout ),
	.cout(Xd_0__inst_inst_add_4_42 ),
	.shareout(Xd_0__inst_inst_add_4_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_41 (
// Equation(s):
// Xd_0__inst_inst_add_2_41_sumout  = SUM(( !Xd_0__inst_r_sum1_5__10__q  $ (!Xd_0__inst_r_sum1_4__10__q  $ (Xd_0__inst_r_sum1_3__10__q )) ) + ( Xd_0__inst_inst_add_2_39  ) + ( Xd_0__inst_inst_add_2_38  ))
// Xd_0__inst_inst_add_2_42  = CARRY(( !Xd_0__inst_r_sum1_5__10__q  $ (!Xd_0__inst_r_sum1_4__10__q  $ (Xd_0__inst_r_sum1_3__10__q )) ) + ( Xd_0__inst_inst_add_2_39  ) + ( Xd_0__inst_inst_add_2_38  ))
// Xd_0__inst_inst_add_2_43  = SHARE((!Xd_0__inst_r_sum1_5__10__q  & (Xd_0__inst_r_sum1_4__10__q  & Xd_0__inst_r_sum1_3__10__q )) # (Xd_0__inst_r_sum1_5__10__q  & ((Xd_0__inst_r_sum1_3__10__q ) # (Xd_0__inst_r_sum1_4__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__10__q ),
	.datac(!Xd_0__inst_r_sum1_4__10__q ),
	.datad(!Xd_0__inst_r_sum1_3__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_38 ),
	.sharein(Xd_0__inst_inst_add_2_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_41_sumout ),
	.cout(Xd_0__inst_inst_add_2_42 ),
	.shareout(Xd_0__inst_inst_add_2_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_42  = CARRY(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_43  = SHARE((!Xd_0__inst_r_sum1_2__10__q  & (Xd_0__inst_r_sum1_1__10__q  & Xd_0__inst_r_sum1_0__10__q )) # (Xd_0__inst_r_sum1_2__10__q  & ((Xd_0__inst_r_sum1_0__10__q ) # (Xd_0__inst_r_sum1_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__10__q ),
	.datac(!Xd_0__inst_r_sum1_1__10__q ),
	.datad(!Xd_0__inst_r_sum1_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_45 (
// Equation(s):
// Xd_0__inst_inst_add_4_45_sumout  = SUM(( !Xd_0__inst_r_sum1_6__11__q  $ (!Xd_0__inst_r_sum1_7__11__q ) ) + ( Xd_0__inst_inst_add_4_43  ) + ( Xd_0__inst_inst_add_4_42  ))
// Xd_0__inst_inst_add_4_46  = CARRY(( !Xd_0__inst_r_sum1_6__11__q  $ (!Xd_0__inst_r_sum1_7__11__q ) ) + ( Xd_0__inst_inst_add_4_43  ) + ( Xd_0__inst_inst_add_4_42  ))
// Xd_0__inst_inst_add_4_47  = SHARE((Xd_0__inst_r_sum1_6__11__q  & Xd_0__inst_r_sum1_7__11__q ))

	.dataa(!Xd_0__inst_r_sum1_6__11__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_42 ),
	.sharein(Xd_0__inst_inst_add_4_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_45_sumout ),
	.cout(Xd_0__inst_inst_add_4_46 ),
	.shareout(Xd_0__inst_inst_add_4_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_45 (
// Equation(s):
// Xd_0__inst_inst_add_2_45_sumout  = SUM(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_43  ) + ( Xd_0__inst_inst_add_2_42  ))
// Xd_0__inst_inst_add_2_46  = CARRY(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_43  ) + ( Xd_0__inst_inst_add_2_42  ))
// Xd_0__inst_inst_add_2_47  = SHARE((!Xd_0__inst_r_sum1_5__11__q  & (Xd_0__inst_r_sum1_4__11__q  & Xd_0__inst_r_sum1_3__11__q )) # (Xd_0__inst_r_sum1_5__11__q  & ((Xd_0__inst_r_sum1_3__11__q ) # (Xd_0__inst_r_sum1_4__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__11__q ),
	.datad(!Xd_0__inst_r_sum1_3__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_42 ),
	.sharein(Xd_0__inst_inst_add_2_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_45_sumout ),
	.cout(Xd_0__inst_inst_add_2_46 ),
	.shareout(Xd_0__inst_inst_add_2_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_46  = CARRY(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_47  = SHARE((!Xd_0__inst_r_sum1_2__11__q  & (Xd_0__inst_r_sum1_1__11__q  & Xd_0__inst_r_sum1_0__11__q )) # (Xd_0__inst_r_sum1_2__11__q  & ((Xd_0__inst_r_sum1_0__11__q ) # (Xd_0__inst_r_sum1_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__11__q ),
	.datad(!Xd_0__inst_r_sum1_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_49 (
// Equation(s):
// Xd_0__inst_inst_add_4_49_sumout  = SUM(( !Xd_0__inst_r_sum1_6__12__q  $ (!Xd_0__inst_r_sum1_7__12__q ) ) + ( Xd_0__inst_inst_add_4_47  ) + ( Xd_0__inst_inst_add_4_46  ))
// Xd_0__inst_inst_add_4_50  = CARRY(( !Xd_0__inst_r_sum1_6__12__q  $ (!Xd_0__inst_r_sum1_7__12__q ) ) + ( Xd_0__inst_inst_add_4_47  ) + ( Xd_0__inst_inst_add_4_46  ))
// Xd_0__inst_inst_add_4_51  = SHARE((Xd_0__inst_r_sum1_6__12__q  & Xd_0__inst_r_sum1_7__12__q ))

	.dataa(!Xd_0__inst_r_sum1_6__12__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_46 ),
	.sharein(Xd_0__inst_inst_add_4_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_49_sumout ),
	.cout(Xd_0__inst_inst_add_4_50 ),
	.shareout(Xd_0__inst_inst_add_4_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_49 (
// Equation(s):
// Xd_0__inst_inst_add_2_49_sumout  = SUM(( !Xd_0__inst_r_sum1_5__12__q  $ (!Xd_0__inst_r_sum1_4__12__q  $ (Xd_0__inst_r_sum1_3__12__q )) ) + ( Xd_0__inst_inst_add_2_47  ) + ( Xd_0__inst_inst_add_2_46  ))
// Xd_0__inst_inst_add_2_50  = CARRY(( !Xd_0__inst_r_sum1_5__12__q  $ (!Xd_0__inst_r_sum1_4__12__q  $ (Xd_0__inst_r_sum1_3__12__q )) ) + ( Xd_0__inst_inst_add_2_47  ) + ( Xd_0__inst_inst_add_2_46  ))
// Xd_0__inst_inst_add_2_51  = SHARE((!Xd_0__inst_r_sum1_5__12__q  & (Xd_0__inst_r_sum1_4__12__q  & Xd_0__inst_r_sum1_3__12__q )) # (Xd_0__inst_r_sum1_5__12__q  & ((Xd_0__inst_r_sum1_3__12__q ) # (Xd_0__inst_r_sum1_4__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__12__q ),
	.datac(!Xd_0__inst_r_sum1_4__12__q ),
	.datad(!Xd_0__inst_r_sum1_3__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_46 ),
	.sharein(Xd_0__inst_inst_add_2_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_49_sumout ),
	.cout(Xd_0__inst_inst_add_2_50 ),
	.shareout(Xd_0__inst_inst_add_2_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_r_sum1_2__12__q  $ (!Xd_0__inst_r_sum1_1__12__q  $ (Xd_0__inst_r_sum1_0__12__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_50  = CARRY(( !Xd_0__inst_r_sum1_2__12__q  $ (!Xd_0__inst_r_sum1_1__12__q  $ (Xd_0__inst_r_sum1_0__12__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_51  = SHARE((!Xd_0__inst_r_sum1_2__12__q  & (Xd_0__inst_r_sum1_1__12__q  & Xd_0__inst_r_sum1_0__12__q )) # (Xd_0__inst_r_sum1_2__12__q  & ((Xd_0__inst_r_sum1_0__12__q ) # (Xd_0__inst_r_sum1_1__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__12__q ),
	.datac(!Xd_0__inst_r_sum1_1__12__q ),
	.datad(!Xd_0__inst_r_sum1_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_53 (
// Equation(s):
// Xd_0__inst_inst_add_4_53_sumout  = SUM(( !Xd_0__inst_r_sum1_6__13__q  $ (!Xd_0__inst_r_sum1_7__13__q ) ) + ( Xd_0__inst_inst_add_4_51  ) + ( Xd_0__inst_inst_add_4_50  ))
// Xd_0__inst_inst_add_4_54  = CARRY(( !Xd_0__inst_r_sum1_6__13__q  $ (!Xd_0__inst_r_sum1_7__13__q ) ) + ( Xd_0__inst_inst_add_4_51  ) + ( Xd_0__inst_inst_add_4_50  ))
// Xd_0__inst_inst_add_4_55  = SHARE((Xd_0__inst_r_sum1_6__13__q  & Xd_0__inst_r_sum1_7__13__q ))

	.dataa(!Xd_0__inst_r_sum1_6__13__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_50 ),
	.sharein(Xd_0__inst_inst_add_4_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_53_sumout ),
	.cout(Xd_0__inst_inst_add_4_54 ),
	.shareout(Xd_0__inst_inst_add_4_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_53 (
// Equation(s):
// Xd_0__inst_inst_add_2_53_sumout  = SUM(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_51  ) + ( Xd_0__inst_inst_add_2_50  ))
// Xd_0__inst_inst_add_2_54  = CARRY(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_51  ) + ( Xd_0__inst_inst_add_2_50  ))
// Xd_0__inst_inst_add_2_55  = SHARE((!Xd_0__inst_r_sum1_5__13__q  & (Xd_0__inst_r_sum1_4__13__q  & Xd_0__inst_r_sum1_3__13__q )) # (Xd_0__inst_r_sum1_5__13__q  & ((Xd_0__inst_r_sum1_3__13__q ) # (Xd_0__inst_r_sum1_4__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__13__q ),
	.datac(!Xd_0__inst_r_sum1_4__13__q ),
	.datad(!Xd_0__inst_r_sum1_3__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_50 ),
	.sharein(Xd_0__inst_inst_add_2_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_53_sumout ),
	.cout(Xd_0__inst_inst_add_2_54 ),
	.shareout(Xd_0__inst_inst_add_2_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))
// Xd_0__inst_inst_add_0_54  = CARRY(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))
// Xd_0__inst_inst_add_0_55  = SHARE((!Xd_0__inst_r_sum1_2__13__q  & (Xd_0__inst_r_sum1_1__13__q  & Xd_0__inst_r_sum1_0__13__q )) # (Xd_0__inst_r_sum1_2__13__q  & ((Xd_0__inst_r_sum1_0__13__q ) # (Xd_0__inst_r_sum1_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__13__q ),
	.datad(!Xd_0__inst_r_sum1_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_57 (
// Equation(s):
// Xd_0__inst_inst_add_4_57_sumout  = SUM(( !Xd_0__inst_r_sum1_6__14__q  $ (!Xd_0__inst_r_sum1_7__14__q ) ) + ( Xd_0__inst_inst_add_4_55  ) + ( Xd_0__inst_inst_add_4_54  ))
// Xd_0__inst_inst_add_4_58  = CARRY(( !Xd_0__inst_r_sum1_6__14__q  $ (!Xd_0__inst_r_sum1_7__14__q ) ) + ( Xd_0__inst_inst_add_4_55  ) + ( Xd_0__inst_inst_add_4_54  ))
// Xd_0__inst_inst_add_4_59  = SHARE((Xd_0__inst_r_sum1_6__14__q  & Xd_0__inst_r_sum1_7__14__q ))

	.dataa(!Xd_0__inst_r_sum1_6__14__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_54 ),
	.sharein(Xd_0__inst_inst_add_4_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_57_sumout ),
	.cout(Xd_0__inst_inst_add_4_58 ),
	.shareout(Xd_0__inst_inst_add_4_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_57 (
// Equation(s):
// Xd_0__inst_inst_add_2_57_sumout  = SUM(( !Xd_0__inst_r_sum1_5__14__q  $ (!Xd_0__inst_r_sum1_4__14__q  $ (Xd_0__inst_r_sum1_3__14__q )) ) + ( Xd_0__inst_inst_add_2_55  ) + ( Xd_0__inst_inst_add_2_54  ))
// Xd_0__inst_inst_add_2_58  = CARRY(( !Xd_0__inst_r_sum1_5__14__q  $ (!Xd_0__inst_r_sum1_4__14__q  $ (Xd_0__inst_r_sum1_3__14__q )) ) + ( Xd_0__inst_inst_add_2_55  ) + ( Xd_0__inst_inst_add_2_54  ))
// Xd_0__inst_inst_add_2_59  = SHARE((!Xd_0__inst_r_sum1_5__14__q  & (Xd_0__inst_r_sum1_4__14__q  & Xd_0__inst_r_sum1_3__14__q )) # (Xd_0__inst_r_sum1_5__14__q  & ((Xd_0__inst_r_sum1_3__14__q ) # (Xd_0__inst_r_sum1_4__14__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__14__q ),
	.datac(!Xd_0__inst_r_sum1_4__14__q ),
	.datad(!Xd_0__inst_r_sum1_3__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_54 ),
	.sharein(Xd_0__inst_inst_add_2_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_57_sumout ),
	.cout(Xd_0__inst_inst_add_2_58 ),
	.shareout(Xd_0__inst_inst_add_2_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_r_sum1_2__14__q  $ (!Xd_0__inst_r_sum1_1__14__q  $ (Xd_0__inst_r_sum1_0__14__q )) ) + ( Xd_0__inst_inst_add_0_55  ) + ( Xd_0__inst_inst_add_0_54  ))
// Xd_0__inst_inst_add_0_58  = CARRY(( !Xd_0__inst_r_sum1_2__14__q  $ (!Xd_0__inst_r_sum1_1__14__q  $ (Xd_0__inst_r_sum1_0__14__q )) ) + ( Xd_0__inst_inst_add_0_55  ) + ( Xd_0__inst_inst_add_0_54  ))
// Xd_0__inst_inst_add_0_59  = SHARE((!Xd_0__inst_r_sum1_2__14__q  & (Xd_0__inst_r_sum1_1__14__q  & Xd_0__inst_r_sum1_0__14__q )) # (Xd_0__inst_r_sum1_2__14__q  & ((Xd_0__inst_r_sum1_0__14__q ) # (Xd_0__inst_r_sum1_1__14__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__14__q ),
	.datac(!Xd_0__inst_r_sum1_1__14__q ),
	.datad(!Xd_0__inst_r_sum1_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_61 (
// Equation(s):
// Xd_0__inst_inst_add_4_61_sumout  = SUM(( !Xd_0__inst_r_sum1_6__15__q  $ (!Xd_0__inst_r_sum1_7__15__q ) ) + ( Xd_0__inst_inst_add_4_59  ) + ( Xd_0__inst_inst_add_4_58  ))
// Xd_0__inst_inst_add_4_62  = CARRY(( !Xd_0__inst_r_sum1_6__15__q  $ (!Xd_0__inst_r_sum1_7__15__q ) ) + ( Xd_0__inst_inst_add_4_59  ) + ( Xd_0__inst_inst_add_4_58  ))
// Xd_0__inst_inst_add_4_63  = SHARE((Xd_0__inst_r_sum1_6__15__q  & Xd_0__inst_r_sum1_7__15__q ))

	.dataa(!Xd_0__inst_r_sum1_6__15__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_58 ),
	.sharein(Xd_0__inst_inst_add_4_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_61_sumout ),
	.cout(Xd_0__inst_inst_add_4_62 ),
	.shareout(Xd_0__inst_inst_add_4_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_61 (
// Equation(s):
// Xd_0__inst_inst_add_2_61_sumout  = SUM(( !Xd_0__inst_r_sum1_5__15__q  $ (!Xd_0__inst_r_sum1_4__15__q  $ (Xd_0__inst_r_sum1_3__15__q )) ) + ( Xd_0__inst_inst_add_2_59  ) + ( Xd_0__inst_inst_add_2_58  ))
// Xd_0__inst_inst_add_2_62  = CARRY(( !Xd_0__inst_r_sum1_5__15__q  $ (!Xd_0__inst_r_sum1_4__15__q  $ (Xd_0__inst_r_sum1_3__15__q )) ) + ( Xd_0__inst_inst_add_2_59  ) + ( Xd_0__inst_inst_add_2_58  ))
// Xd_0__inst_inst_add_2_63  = SHARE((!Xd_0__inst_r_sum1_5__15__q  & (Xd_0__inst_r_sum1_4__15__q  & Xd_0__inst_r_sum1_3__15__q )) # (Xd_0__inst_r_sum1_5__15__q  & ((Xd_0__inst_r_sum1_3__15__q ) # (Xd_0__inst_r_sum1_4__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__15__q ),
	.datac(!Xd_0__inst_r_sum1_4__15__q ),
	.datad(!Xd_0__inst_r_sum1_3__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_58 ),
	.sharein(Xd_0__inst_inst_add_2_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_61_sumout ),
	.cout(Xd_0__inst_inst_add_2_62 ),
	.shareout(Xd_0__inst_inst_add_2_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_r_sum1_2__15__q  $ (!Xd_0__inst_r_sum1_1__15__q  $ (Xd_0__inst_r_sum1_0__15__q )) ) + ( Xd_0__inst_inst_add_0_59  ) + ( Xd_0__inst_inst_add_0_58  ))
// Xd_0__inst_inst_add_0_62  = CARRY(( !Xd_0__inst_r_sum1_2__15__q  $ (!Xd_0__inst_r_sum1_1__15__q  $ (Xd_0__inst_r_sum1_0__15__q )) ) + ( Xd_0__inst_inst_add_0_59  ) + ( Xd_0__inst_inst_add_0_58  ))
// Xd_0__inst_inst_add_0_63  = SHARE((!Xd_0__inst_r_sum1_2__15__q  & (Xd_0__inst_r_sum1_1__15__q  & Xd_0__inst_r_sum1_0__15__q )) # (Xd_0__inst_r_sum1_2__15__q  & ((Xd_0__inst_r_sum1_0__15__q ) # (Xd_0__inst_r_sum1_1__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__15__q ),
	.datac(!Xd_0__inst_r_sum1_1__15__q ),
	.datad(!Xd_0__inst_r_sum1_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_add_0_62 ),
	.shareout(Xd_0__inst_inst_add_0_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_65 (
// Equation(s):
// Xd_0__inst_inst_add_4_65_sumout  = SUM(( !Xd_0__inst_r_sum1_6__16__q  $ (!Xd_0__inst_r_sum1_7__16__q ) ) + ( Xd_0__inst_inst_add_4_63  ) + ( Xd_0__inst_inst_add_4_62  ))
// Xd_0__inst_inst_add_4_66  = CARRY(( !Xd_0__inst_r_sum1_6__16__q  $ (!Xd_0__inst_r_sum1_7__16__q ) ) + ( Xd_0__inst_inst_add_4_63  ) + ( Xd_0__inst_inst_add_4_62  ))
// Xd_0__inst_inst_add_4_67  = SHARE((Xd_0__inst_r_sum1_6__16__q  & Xd_0__inst_r_sum1_7__16__q ))

	.dataa(!Xd_0__inst_r_sum1_6__16__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_62 ),
	.sharein(Xd_0__inst_inst_add_4_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_65_sumout ),
	.cout(Xd_0__inst_inst_add_4_66 ),
	.shareout(Xd_0__inst_inst_add_4_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_65 (
// Equation(s):
// Xd_0__inst_inst_add_2_65_sumout  = SUM(( !Xd_0__inst_r_sum1_5__16__q  $ (!Xd_0__inst_r_sum1_4__16__q  $ (Xd_0__inst_r_sum1_3__16__q )) ) + ( Xd_0__inst_inst_add_2_63  ) + ( Xd_0__inst_inst_add_2_62  ))
// Xd_0__inst_inst_add_2_66  = CARRY(( !Xd_0__inst_r_sum1_5__16__q  $ (!Xd_0__inst_r_sum1_4__16__q  $ (Xd_0__inst_r_sum1_3__16__q )) ) + ( Xd_0__inst_inst_add_2_63  ) + ( Xd_0__inst_inst_add_2_62  ))
// Xd_0__inst_inst_add_2_67  = SHARE((!Xd_0__inst_r_sum1_5__16__q  & (Xd_0__inst_r_sum1_4__16__q  & Xd_0__inst_r_sum1_3__16__q )) # (Xd_0__inst_r_sum1_5__16__q  & ((Xd_0__inst_r_sum1_3__16__q ) # (Xd_0__inst_r_sum1_4__16__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__16__q ),
	.datac(!Xd_0__inst_r_sum1_4__16__q ),
	.datad(!Xd_0__inst_r_sum1_3__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_62 ),
	.sharein(Xd_0__inst_inst_add_2_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_65_sumout ),
	.cout(Xd_0__inst_inst_add_2_66 ),
	.shareout(Xd_0__inst_inst_add_2_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_65 (
// Equation(s):
// Xd_0__inst_inst_add_0_65_sumout  = SUM(( !Xd_0__inst_r_sum1_2__16__q  $ (!Xd_0__inst_r_sum1_1__16__q  $ (Xd_0__inst_r_sum1_0__16__q )) ) + ( Xd_0__inst_inst_add_0_63  ) + ( Xd_0__inst_inst_add_0_62  ))
// Xd_0__inst_inst_add_0_66  = CARRY(( !Xd_0__inst_r_sum1_2__16__q  $ (!Xd_0__inst_r_sum1_1__16__q  $ (Xd_0__inst_r_sum1_0__16__q )) ) + ( Xd_0__inst_inst_add_0_63  ) + ( Xd_0__inst_inst_add_0_62  ))
// Xd_0__inst_inst_add_0_67  = SHARE((!Xd_0__inst_r_sum1_2__16__q  & (Xd_0__inst_r_sum1_1__16__q  & Xd_0__inst_r_sum1_0__16__q )) # (Xd_0__inst_r_sum1_2__16__q  & ((Xd_0__inst_r_sum1_0__16__q ) # (Xd_0__inst_r_sum1_1__16__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__16__q ),
	.datac(!Xd_0__inst_r_sum1_1__16__q ),
	.datad(!Xd_0__inst_r_sum1_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_62 ),
	.sharein(Xd_0__inst_inst_add_0_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_65_sumout ),
	.cout(Xd_0__inst_inst_add_0_66 ),
	.shareout(Xd_0__inst_inst_add_0_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_69 (
// Equation(s):
// Xd_0__inst_inst_add_4_69_sumout  = SUM(( !Xd_0__inst_r_sum1_6__17__q  $ (!Xd_0__inst_r_sum1_7__17__q ) ) + ( Xd_0__inst_inst_add_4_67  ) + ( Xd_0__inst_inst_add_4_66  ))
// Xd_0__inst_inst_add_4_70  = CARRY(( !Xd_0__inst_r_sum1_6__17__q  $ (!Xd_0__inst_r_sum1_7__17__q ) ) + ( Xd_0__inst_inst_add_4_67  ) + ( Xd_0__inst_inst_add_4_66  ))
// Xd_0__inst_inst_add_4_71  = SHARE((Xd_0__inst_r_sum1_6__17__q  & Xd_0__inst_r_sum1_7__17__q ))

	.dataa(!Xd_0__inst_r_sum1_6__17__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_66 ),
	.sharein(Xd_0__inst_inst_add_4_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_69_sumout ),
	.cout(Xd_0__inst_inst_add_4_70 ),
	.shareout(Xd_0__inst_inst_add_4_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_69 (
// Equation(s):
// Xd_0__inst_inst_add_2_69_sumout  = SUM(( !Xd_0__inst_r_sum1_5__17__q  $ (!Xd_0__inst_r_sum1_4__17__q  $ (Xd_0__inst_r_sum1_3__17__q )) ) + ( Xd_0__inst_inst_add_2_67  ) + ( Xd_0__inst_inst_add_2_66  ))
// Xd_0__inst_inst_add_2_70  = CARRY(( !Xd_0__inst_r_sum1_5__17__q  $ (!Xd_0__inst_r_sum1_4__17__q  $ (Xd_0__inst_r_sum1_3__17__q )) ) + ( Xd_0__inst_inst_add_2_67  ) + ( Xd_0__inst_inst_add_2_66  ))
// Xd_0__inst_inst_add_2_71  = SHARE((!Xd_0__inst_r_sum1_5__17__q  & (Xd_0__inst_r_sum1_4__17__q  & Xd_0__inst_r_sum1_3__17__q )) # (Xd_0__inst_r_sum1_5__17__q  & ((Xd_0__inst_r_sum1_3__17__q ) # (Xd_0__inst_r_sum1_4__17__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__17__q ),
	.datac(!Xd_0__inst_r_sum1_4__17__q ),
	.datad(!Xd_0__inst_r_sum1_3__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_66 ),
	.sharein(Xd_0__inst_inst_add_2_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_69_sumout ),
	.cout(Xd_0__inst_inst_add_2_70 ),
	.shareout(Xd_0__inst_inst_add_2_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_69 (
// Equation(s):
// Xd_0__inst_inst_add_0_69_sumout  = SUM(( !Xd_0__inst_r_sum1_2__17__q  $ (!Xd_0__inst_r_sum1_1__17__q  $ (Xd_0__inst_r_sum1_0__17__q )) ) + ( Xd_0__inst_inst_add_0_67  ) + ( Xd_0__inst_inst_add_0_66  ))
// Xd_0__inst_inst_add_0_70  = CARRY(( !Xd_0__inst_r_sum1_2__17__q  $ (!Xd_0__inst_r_sum1_1__17__q  $ (Xd_0__inst_r_sum1_0__17__q )) ) + ( Xd_0__inst_inst_add_0_67  ) + ( Xd_0__inst_inst_add_0_66  ))
// Xd_0__inst_inst_add_0_71  = SHARE((!Xd_0__inst_r_sum1_2__17__q  & (Xd_0__inst_r_sum1_1__17__q  & Xd_0__inst_r_sum1_0__17__q )) # (Xd_0__inst_r_sum1_2__17__q  & ((Xd_0__inst_r_sum1_0__17__q ) # (Xd_0__inst_r_sum1_1__17__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__17__q ),
	.datac(!Xd_0__inst_r_sum1_1__17__q ),
	.datad(!Xd_0__inst_r_sum1_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_66 ),
	.sharein(Xd_0__inst_inst_add_0_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_69_sumout ),
	.cout(Xd_0__inst_inst_add_0_70 ),
	.shareout(Xd_0__inst_inst_add_0_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_73 (
// Equation(s):
// Xd_0__inst_inst_add_4_73_sumout  = SUM(( !Xd_0__inst_r_sum1_6__18__q  $ (!Xd_0__inst_r_sum1_7__18__q ) ) + ( Xd_0__inst_inst_add_4_71  ) + ( Xd_0__inst_inst_add_4_70  ))
// Xd_0__inst_inst_add_4_74  = CARRY(( !Xd_0__inst_r_sum1_6__18__q  $ (!Xd_0__inst_r_sum1_7__18__q ) ) + ( Xd_0__inst_inst_add_4_71  ) + ( Xd_0__inst_inst_add_4_70  ))
// Xd_0__inst_inst_add_4_75  = SHARE((Xd_0__inst_r_sum1_6__18__q  & Xd_0__inst_r_sum1_7__18__q ))

	.dataa(!Xd_0__inst_r_sum1_6__18__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_70 ),
	.sharein(Xd_0__inst_inst_add_4_71 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_73_sumout ),
	.cout(Xd_0__inst_inst_add_4_74 ),
	.shareout(Xd_0__inst_inst_add_4_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_73 (
// Equation(s):
// Xd_0__inst_inst_add_2_73_sumout  = SUM(( !Xd_0__inst_r_sum1_5__18__q  $ (!Xd_0__inst_r_sum1_4__18__q  $ (Xd_0__inst_r_sum1_3__18__q )) ) + ( Xd_0__inst_inst_add_2_71  ) + ( Xd_0__inst_inst_add_2_70  ))
// Xd_0__inst_inst_add_2_74  = CARRY(( !Xd_0__inst_r_sum1_5__18__q  $ (!Xd_0__inst_r_sum1_4__18__q  $ (Xd_0__inst_r_sum1_3__18__q )) ) + ( Xd_0__inst_inst_add_2_71  ) + ( Xd_0__inst_inst_add_2_70  ))
// Xd_0__inst_inst_add_2_75  = SHARE((!Xd_0__inst_r_sum1_5__18__q  & (Xd_0__inst_r_sum1_4__18__q  & Xd_0__inst_r_sum1_3__18__q )) # (Xd_0__inst_r_sum1_5__18__q  & ((Xd_0__inst_r_sum1_3__18__q ) # (Xd_0__inst_r_sum1_4__18__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__18__q ),
	.datac(!Xd_0__inst_r_sum1_4__18__q ),
	.datad(!Xd_0__inst_r_sum1_3__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_70 ),
	.sharein(Xd_0__inst_inst_add_2_71 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_73_sumout ),
	.cout(Xd_0__inst_inst_add_2_74 ),
	.shareout(Xd_0__inst_inst_add_2_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_73 (
// Equation(s):
// Xd_0__inst_inst_add_0_73_sumout  = SUM(( !Xd_0__inst_r_sum1_2__18__q  $ (!Xd_0__inst_r_sum1_1__18__q  $ (Xd_0__inst_r_sum1_0__18__q )) ) + ( Xd_0__inst_inst_add_0_71  ) + ( Xd_0__inst_inst_add_0_70  ))
// Xd_0__inst_inst_add_0_74  = CARRY(( !Xd_0__inst_r_sum1_2__18__q  $ (!Xd_0__inst_r_sum1_1__18__q  $ (Xd_0__inst_r_sum1_0__18__q )) ) + ( Xd_0__inst_inst_add_0_71  ) + ( Xd_0__inst_inst_add_0_70  ))
// Xd_0__inst_inst_add_0_75  = SHARE((!Xd_0__inst_r_sum1_2__18__q  & (Xd_0__inst_r_sum1_1__18__q  & Xd_0__inst_r_sum1_0__18__q )) # (Xd_0__inst_r_sum1_2__18__q  & ((Xd_0__inst_r_sum1_0__18__q ) # (Xd_0__inst_r_sum1_1__18__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__18__q ),
	.datac(!Xd_0__inst_r_sum1_1__18__q ),
	.datad(!Xd_0__inst_r_sum1_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_70 ),
	.sharein(Xd_0__inst_inst_add_0_71 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_73_sumout ),
	.cout(Xd_0__inst_inst_add_0_74 ),
	.shareout(Xd_0__inst_inst_add_0_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_77 (
// Equation(s):
// Xd_0__inst_inst_add_4_77_sumout  = SUM(( !Xd_0__inst_r_sum1_6__19__q  $ (!Xd_0__inst_r_sum1_7__19__q ) ) + ( Xd_0__inst_inst_add_4_75  ) + ( Xd_0__inst_inst_add_4_74  ))
// Xd_0__inst_inst_add_4_78  = CARRY(( !Xd_0__inst_r_sum1_6__19__q  $ (!Xd_0__inst_r_sum1_7__19__q ) ) + ( Xd_0__inst_inst_add_4_75  ) + ( Xd_0__inst_inst_add_4_74  ))
// Xd_0__inst_inst_add_4_79  = SHARE((Xd_0__inst_r_sum1_6__19__q  & Xd_0__inst_r_sum1_7__19__q ))

	.dataa(!Xd_0__inst_r_sum1_6__19__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_74 ),
	.sharein(Xd_0__inst_inst_add_4_75 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_77_sumout ),
	.cout(Xd_0__inst_inst_add_4_78 ),
	.shareout(Xd_0__inst_inst_add_4_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_77 (
// Equation(s):
// Xd_0__inst_inst_add_2_77_sumout  = SUM(( !Xd_0__inst_r_sum1_5__19__q  $ (!Xd_0__inst_r_sum1_4__19__q  $ (Xd_0__inst_r_sum1_3__19__q )) ) + ( Xd_0__inst_inst_add_2_75  ) + ( Xd_0__inst_inst_add_2_74  ))
// Xd_0__inst_inst_add_2_78  = CARRY(( !Xd_0__inst_r_sum1_5__19__q  $ (!Xd_0__inst_r_sum1_4__19__q  $ (Xd_0__inst_r_sum1_3__19__q )) ) + ( Xd_0__inst_inst_add_2_75  ) + ( Xd_0__inst_inst_add_2_74  ))
// Xd_0__inst_inst_add_2_79  = SHARE((!Xd_0__inst_r_sum1_5__19__q  & (Xd_0__inst_r_sum1_4__19__q  & Xd_0__inst_r_sum1_3__19__q )) # (Xd_0__inst_r_sum1_5__19__q  & ((Xd_0__inst_r_sum1_3__19__q ) # (Xd_0__inst_r_sum1_4__19__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__19__q ),
	.datac(!Xd_0__inst_r_sum1_4__19__q ),
	.datad(!Xd_0__inst_r_sum1_3__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_74 ),
	.sharein(Xd_0__inst_inst_add_2_75 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_77_sumout ),
	.cout(Xd_0__inst_inst_add_2_78 ),
	.shareout(Xd_0__inst_inst_add_2_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_77 (
// Equation(s):
// Xd_0__inst_inst_add_0_77_sumout  = SUM(( !Xd_0__inst_r_sum1_2__19__q  $ (!Xd_0__inst_r_sum1_1__19__q  $ (Xd_0__inst_r_sum1_0__19__q )) ) + ( Xd_0__inst_inst_add_0_75  ) + ( Xd_0__inst_inst_add_0_74  ))
// Xd_0__inst_inst_add_0_78  = CARRY(( !Xd_0__inst_r_sum1_2__19__q  $ (!Xd_0__inst_r_sum1_1__19__q  $ (Xd_0__inst_r_sum1_0__19__q )) ) + ( Xd_0__inst_inst_add_0_75  ) + ( Xd_0__inst_inst_add_0_74  ))
// Xd_0__inst_inst_add_0_79  = SHARE((!Xd_0__inst_r_sum1_2__19__q  & (Xd_0__inst_r_sum1_1__19__q  & Xd_0__inst_r_sum1_0__19__q )) # (Xd_0__inst_r_sum1_2__19__q  & ((Xd_0__inst_r_sum1_0__19__q ) # (Xd_0__inst_r_sum1_1__19__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__19__q ),
	.datac(!Xd_0__inst_r_sum1_1__19__q ),
	.datad(!Xd_0__inst_r_sum1_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_74 ),
	.sharein(Xd_0__inst_inst_add_0_75 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_77_sumout ),
	.cout(Xd_0__inst_inst_add_0_78 ),
	.shareout(Xd_0__inst_inst_add_0_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_81 (
// Equation(s):
// Xd_0__inst_inst_add_4_81_sumout  = SUM(( !Xd_0__inst_r_sum1_6__20__q  $ (!Xd_0__inst_r_sum1_7__20__q ) ) + ( Xd_0__inst_inst_add_4_79  ) + ( Xd_0__inst_inst_add_4_78  ))
// Xd_0__inst_inst_add_4_82  = CARRY(( !Xd_0__inst_r_sum1_6__20__q  $ (!Xd_0__inst_r_sum1_7__20__q ) ) + ( Xd_0__inst_inst_add_4_79  ) + ( Xd_0__inst_inst_add_4_78  ))
// Xd_0__inst_inst_add_4_83  = SHARE((Xd_0__inst_r_sum1_6__20__q  & Xd_0__inst_r_sum1_7__20__q ))

	.dataa(!Xd_0__inst_r_sum1_6__20__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_78 ),
	.sharein(Xd_0__inst_inst_add_4_79 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_81_sumout ),
	.cout(Xd_0__inst_inst_add_4_82 ),
	.shareout(Xd_0__inst_inst_add_4_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_81 (
// Equation(s):
// Xd_0__inst_inst_add_2_81_sumout  = SUM(( !Xd_0__inst_r_sum1_5__20__q  $ (!Xd_0__inst_r_sum1_4__20__q  $ (Xd_0__inst_r_sum1_3__20__q )) ) + ( Xd_0__inst_inst_add_2_79  ) + ( Xd_0__inst_inst_add_2_78  ))
// Xd_0__inst_inst_add_2_82  = CARRY(( !Xd_0__inst_r_sum1_5__20__q  $ (!Xd_0__inst_r_sum1_4__20__q  $ (Xd_0__inst_r_sum1_3__20__q )) ) + ( Xd_0__inst_inst_add_2_79  ) + ( Xd_0__inst_inst_add_2_78  ))
// Xd_0__inst_inst_add_2_83  = SHARE((!Xd_0__inst_r_sum1_5__20__q  & (Xd_0__inst_r_sum1_4__20__q  & Xd_0__inst_r_sum1_3__20__q )) # (Xd_0__inst_r_sum1_5__20__q  & ((Xd_0__inst_r_sum1_3__20__q ) # (Xd_0__inst_r_sum1_4__20__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__20__q ),
	.datac(!Xd_0__inst_r_sum1_4__20__q ),
	.datad(!Xd_0__inst_r_sum1_3__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_78 ),
	.sharein(Xd_0__inst_inst_add_2_79 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_81_sumout ),
	.cout(Xd_0__inst_inst_add_2_82 ),
	.shareout(Xd_0__inst_inst_add_2_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_81 (
// Equation(s):
// Xd_0__inst_inst_add_0_81_sumout  = SUM(( !Xd_0__inst_r_sum1_2__20__q  $ (!Xd_0__inst_r_sum1_1__20__q  $ (Xd_0__inst_r_sum1_0__20__q )) ) + ( Xd_0__inst_inst_add_0_79  ) + ( Xd_0__inst_inst_add_0_78  ))
// Xd_0__inst_inst_add_0_82  = CARRY(( !Xd_0__inst_r_sum1_2__20__q  $ (!Xd_0__inst_r_sum1_1__20__q  $ (Xd_0__inst_r_sum1_0__20__q )) ) + ( Xd_0__inst_inst_add_0_79  ) + ( Xd_0__inst_inst_add_0_78  ))
// Xd_0__inst_inst_add_0_83  = SHARE((!Xd_0__inst_r_sum1_2__20__q  & (Xd_0__inst_r_sum1_1__20__q  & Xd_0__inst_r_sum1_0__20__q )) # (Xd_0__inst_r_sum1_2__20__q  & ((Xd_0__inst_r_sum1_0__20__q ) # (Xd_0__inst_r_sum1_1__20__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__20__q ),
	.datac(!Xd_0__inst_r_sum1_1__20__q ),
	.datad(!Xd_0__inst_r_sum1_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_78 ),
	.sharein(Xd_0__inst_inst_add_0_79 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_add_0_82 ),
	.shareout(Xd_0__inst_inst_add_0_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_85 (
// Equation(s):
// Xd_0__inst_inst_add_4_85_sumout  = SUM(( !Xd_0__inst_r_sum1_6__21__q  $ (!Xd_0__inst_r_sum1_7__21__q ) ) + ( Xd_0__inst_inst_add_4_83  ) + ( Xd_0__inst_inst_add_4_82  ))
// Xd_0__inst_inst_add_4_86  = CARRY(( !Xd_0__inst_r_sum1_6__21__q  $ (!Xd_0__inst_r_sum1_7__21__q ) ) + ( Xd_0__inst_inst_add_4_83  ) + ( Xd_0__inst_inst_add_4_82  ))
// Xd_0__inst_inst_add_4_87  = SHARE((Xd_0__inst_r_sum1_6__21__q  & Xd_0__inst_r_sum1_7__21__q ))

	.dataa(!Xd_0__inst_r_sum1_6__21__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_82 ),
	.sharein(Xd_0__inst_inst_add_4_83 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_85_sumout ),
	.cout(Xd_0__inst_inst_add_4_86 ),
	.shareout(Xd_0__inst_inst_add_4_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_85 (
// Equation(s):
// Xd_0__inst_inst_add_2_85_sumout  = SUM(( !Xd_0__inst_r_sum1_5__21__q  $ (!Xd_0__inst_r_sum1_4__21__q  $ (Xd_0__inst_r_sum1_3__21__q )) ) + ( Xd_0__inst_inst_add_2_83  ) + ( Xd_0__inst_inst_add_2_82  ))
// Xd_0__inst_inst_add_2_86  = CARRY(( !Xd_0__inst_r_sum1_5__21__q  $ (!Xd_0__inst_r_sum1_4__21__q  $ (Xd_0__inst_r_sum1_3__21__q )) ) + ( Xd_0__inst_inst_add_2_83  ) + ( Xd_0__inst_inst_add_2_82  ))
// Xd_0__inst_inst_add_2_87  = SHARE((!Xd_0__inst_r_sum1_5__21__q  & (Xd_0__inst_r_sum1_4__21__q  & Xd_0__inst_r_sum1_3__21__q )) # (Xd_0__inst_r_sum1_5__21__q  & ((Xd_0__inst_r_sum1_3__21__q ) # (Xd_0__inst_r_sum1_4__21__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__21__q ),
	.datac(!Xd_0__inst_r_sum1_4__21__q ),
	.datad(!Xd_0__inst_r_sum1_3__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_82 ),
	.sharein(Xd_0__inst_inst_add_2_83 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_85_sumout ),
	.cout(Xd_0__inst_inst_add_2_86 ),
	.shareout(Xd_0__inst_inst_add_2_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_85 (
// Equation(s):
// Xd_0__inst_inst_add_0_85_sumout  = SUM(( !Xd_0__inst_r_sum1_2__21__q  $ (!Xd_0__inst_r_sum1_1__21__q  $ (Xd_0__inst_r_sum1_0__21__q )) ) + ( Xd_0__inst_inst_add_0_83  ) + ( Xd_0__inst_inst_add_0_82  ))
// Xd_0__inst_inst_add_0_86  = CARRY(( !Xd_0__inst_r_sum1_2__21__q  $ (!Xd_0__inst_r_sum1_1__21__q  $ (Xd_0__inst_r_sum1_0__21__q )) ) + ( Xd_0__inst_inst_add_0_83  ) + ( Xd_0__inst_inst_add_0_82  ))
// Xd_0__inst_inst_add_0_87  = SHARE((!Xd_0__inst_r_sum1_2__21__q  & (Xd_0__inst_r_sum1_1__21__q  & Xd_0__inst_r_sum1_0__21__q )) # (Xd_0__inst_r_sum1_2__21__q  & ((Xd_0__inst_r_sum1_0__21__q ) # (Xd_0__inst_r_sum1_1__21__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__21__q ),
	.datac(!Xd_0__inst_r_sum1_1__21__q ),
	.datad(!Xd_0__inst_r_sum1_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_82 ),
	.sharein(Xd_0__inst_inst_add_0_83 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_85_sumout ),
	.cout(Xd_0__inst_inst_add_0_86 ),
	.shareout(Xd_0__inst_inst_add_0_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_89 (
// Equation(s):
// Xd_0__inst_inst_add_4_89_sumout  = SUM(( !Xd_0__inst_r_sum1_6__22__q  $ (!Xd_0__inst_r_sum1_7__22__q ) ) + ( Xd_0__inst_inst_add_4_87  ) + ( Xd_0__inst_inst_add_4_86  ))
// Xd_0__inst_inst_add_4_90  = CARRY(( !Xd_0__inst_r_sum1_6__22__q  $ (!Xd_0__inst_r_sum1_7__22__q ) ) + ( Xd_0__inst_inst_add_4_87  ) + ( Xd_0__inst_inst_add_4_86  ))
// Xd_0__inst_inst_add_4_91  = SHARE((Xd_0__inst_r_sum1_6__22__q  & Xd_0__inst_r_sum1_7__22__q ))

	.dataa(!Xd_0__inst_r_sum1_6__22__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_86 ),
	.sharein(Xd_0__inst_inst_add_4_87 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_89_sumout ),
	.cout(Xd_0__inst_inst_add_4_90 ),
	.shareout(Xd_0__inst_inst_add_4_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_89 (
// Equation(s):
// Xd_0__inst_inst_add_2_89_sumout  = SUM(( !Xd_0__inst_r_sum1_5__22__q  $ (!Xd_0__inst_r_sum1_4__22__q  $ (Xd_0__inst_r_sum1_3__22__q )) ) + ( Xd_0__inst_inst_add_2_87  ) + ( Xd_0__inst_inst_add_2_86  ))
// Xd_0__inst_inst_add_2_90  = CARRY(( !Xd_0__inst_r_sum1_5__22__q  $ (!Xd_0__inst_r_sum1_4__22__q  $ (Xd_0__inst_r_sum1_3__22__q )) ) + ( Xd_0__inst_inst_add_2_87  ) + ( Xd_0__inst_inst_add_2_86  ))
// Xd_0__inst_inst_add_2_91  = SHARE((!Xd_0__inst_r_sum1_5__22__q  & (Xd_0__inst_r_sum1_4__22__q  & Xd_0__inst_r_sum1_3__22__q )) # (Xd_0__inst_r_sum1_5__22__q  & ((Xd_0__inst_r_sum1_3__22__q ) # (Xd_0__inst_r_sum1_4__22__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__22__q ),
	.datac(!Xd_0__inst_r_sum1_4__22__q ),
	.datad(!Xd_0__inst_r_sum1_3__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_86 ),
	.sharein(Xd_0__inst_inst_add_2_87 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_89_sumout ),
	.cout(Xd_0__inst_inst_add_2_90 ),
	.shareout(Xd_0__inst_inst_add_2_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_89 (
// Equation(s):
// Xd_0__inst_inst_add_0_89_sumout  = SUM(( !Xd_0__inst_r_sum1_2__22__q  $ (!Xd_0__inst_r_sum1_1__22__q  $ (Xd_0__inst_r_sum1_0__22__q )) ) + ( Xd_0__inst_inst_add_0_87  ) + ( Xd_0__inst_inst_add_0_86  ))
// Xd_0__inst_inst_add_0_90  = CARRY(( !Xd_0__inst_r_sum1_2__22__q  $ (!Xd_0__inst_r_sum1_1__22__q  $ (Xd_0__inst_r_sum1_0__22__q )) ) + ( Xd_0__inst_inst_add_0_87  ) + ( Xd_0__inst_inst_add_0_86  ))
// Xd_0__inst_inst_add_0_91  = SHARE((!Xd_0__inst_r_sum1_2__22__q  & (Xd_0__inst_r_sum1_1__22__q  & Xd_0__inst_r_sum1_0__22__q )) # (Xd_0__inst_r_sum1_2__22__q  & ((Xd_0__inst_r_sum1_0__22__q ) # (Xd_0__inst_r_sum1_1__22__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__22__q ),
	.datac(!Xd_0__inst_r_sum1_1__22__q ),
	.datad(!Xd_0__inst_r_sum1_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_86 ),
	.sharein(Xd_0__inst_inst_add_0_87 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_89_sumout ),
	.cout(Xd_0__inst_inst_add_0_90 ),
	.shareout(Xd_0__inst_inst_add_0_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_93 (
// Equation(s):
// Xd_0__inst_inst_add_4_93_sumout  = SUM(( !Xd_0__inst_r_sum1_6__23__q  $ (!Xd_0__inst_r_sum1_7__23__q ) ) + ( Xd_0__inst_inst_add_4_91  ) + ( Xd_0__inst_inst_add_4_90  ))
// Xd_0__inst_inst_add_4_94  = CARRY(( !Xd_0__inst_r_sum1_6__23__q  $ (!Xd_0__inst_r_sum1_7__23__q ) ) + ( Xd_0__inst_inst_add_4_91  ) + ( Xd_0__inst_inst_add_4_90  ))
// Xd_0__inst_inst_add_4_95  = SHARE((Xd_0__inst_r_sum1_6__23__q  & Xd_0__inst_r_sum1_7__23__q ))

	.dataa(!Xd_0__inst_r_sum1_6__23__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_90 ),
	.sharein(Xd_0__inst_inst_add_4_91 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_93_sumout ),
	.cout(Xd_0__inst_inst_add_4_94 ),
	.shareout(Xd_0__inst_inst_add_4_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_93 (
// Equation(s):
// Xd_0__inst_inst_add_2_93_sumout  = SUM(( !Xd_0__inst_r_sum1_5__23__q  $ (!Xd_0__inst_r_sum1_4__23__q  $ (Xd_0__inst_r_sum1_3__23__q )) ) + ( Xd_0__inst_inst_add_2_91  ) + ( Xd_0__inst_inst_add_2_90  ))
// Xd_0__inst_inst_add_2_94  = CARRY(( !Xd_0__inst_r_sum1_5__23__q  $ (!Xd_0__inst_r_sum1_4__23__q  $ (Xd_0__inst_r_sum1_3__23__q )) ) + ( Xd_0__inst_inst_add_2_91  ) + ( Xd_0__inst_inst_add_2_90  ))
// Xd_0__inst_inst_add_2_95  = SHARE((!Xd_0__inst_r_sum1_5__23__q  & (Xd_0__inst_r_sum1_4__23__q  & Xd_0__inst_r_sum1_3__23__q )) # (Xd_0__inst_r_sum1_5__23__q  & ((Xd_0__inst_r_sum1_3__23__q ) # (Xd_0__inst_r_sum1_4__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__23__q ),
	.datac(!Xd_0__inst_r_sum1_4__23__q ),
	.datad(!Xd_0__inst_r_sum1_3__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_90 ),
	.sharein(Xd_0__inst_inst_add_2_91 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_93_sumout ),
	.cout(Xd_0__inst_inst_add_2_94 ),
	.shareout(Xd_0__inst_inst_add_2_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_93 (
// Equation(s):
// Xd_0__inst_inst_add_0_93_sumout  = SUM(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_91  ) + ( Xd_0__inst_inst_add_0_90  ))
// Xd_0__inst_inst_add_0_94  = CARRY(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_91  ) + ( Xd_0__inst_inst_add_0_90  ))
// Xd_0__inst_inst_add_0_95  = SHARE((!Xd_0__inst_r_sum1_2__23__q  & (Xd_0__inst_r_sum1_1__23__q  & Xd_0__inst_r_sum1_0__23__q )) # (Xd_0__inst_r_sum1_2__23__q  & ((Xd_0__inst_r_sum1_0__23__q ) # (Xd_0__inst_r_sum1_1__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__23__q ),
	.datad(!Xd_0__inst_r_sum1_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_90 ),
	.sharein(Xd_0__inst_inst_add_0_91 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_93_sumout ),
	.cout(Xd_0__inst_inst_add_0_94 ),
	.shareout(Xd_0__inst_inst_add_0_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_97 (
// Equation(s):
// Xd_0__inst_inst_add_4_97_sumout  = SUM(( !Xd_0__inst_r_sum1_6__23__q  $ (!Xd_0__inst_r_sum1_7__23__q ) ) + ( Xd_0__inst_inst_add_4_95  ) + ( Xd_0__inst_inst_add_4_94  ))

	.dataa(!Xd_0__inst_r_sum1_6__23__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_r_sum1_7__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_94 ),
	.sharein(Xd_0__inst_inst_add_4_95 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_97_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_97 (
// Equation(s):
// Xd_0__inst_inst_add_2_97_sumout  = SUM(( !Xd_0__inst_r_sum1_5__23__q  $ (!Xd_0__inst_r_sum1_4__23__q  $ (Xd_0__inst_r_sum1_3__23__q )) ) + ( Xd_0__inst_inst_add_2_95  ) + ( Xd_0__inst_inst_add_2_94  ))
// Xd_0__inst_inst_add_2_98  = CARRY(( !Xd_0__inst_r_sum1_5__23__q  $ (!Xd_0__inst_r_sum1_4__23__q  $ (Xd_0__inst_r_sum1_3__23__q )) ) + ( Xd_0__inst_inst_add_2_95  ) + ( Xd_0__inst_inst_add_2_94  ))
// Xd_0__inst_inst_add_2_99  = SHARE((!Xd_0__inst_r_sum1_5__23__q  & (Xd_0__inst_r_sum1_4__23__q  & Xd_0__inst_r_sum1_3__23__q )) # (Xd_0__inst_r_sum1_5__23__q  & ((Xd_0__inst_r_sum1_3__23__q ) # (Xd_0__inst_r_sum1_4__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__23__q ),
	.datac(!Xd_0__inst_r_sum1_4__23__q ),
	.datad(!Xd_0__inst_r_sum1_3__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_94 ),
	.sharein(Xd_0__inst_inst_add_2_95 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_97_sumout ),
	.cout(Xd_0__inst_inst_add_2_98 ),
	.shareout(Xd_0__inst_inst_add_2_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_97 (
// Equation(s):
// Xd_0__inst_inst_add_0_97_sumout  = SUM(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_95  ) + ( Xd_0__inst_inst_add_0_94  ))
// Xd_0__inst_inst_add_0_98  = CARRY(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_95  ) + ( Xd_0__inst_inst_add_0_94  ))
// Xd_0__inst_inst_add_0_99  = SHARE((!Xd_0__inst_r_sum1_2__23__q  & (Xd_0__inst_r_sum1_1__23__q  & Xd_0__inst_r_sum1_0__23__q )) # (Xd_0__inst_r_sum1_2__23__q  & ((Xd_0__inst_r_sum1_0__23__q ) # (Xd_0__inst_r_sum1_1__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__23__q ),
	.datad(!Xd_0__inst_r_sum1_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_94 ),
	.sharein(Xd_0__inst_inst_add_0_95 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_97_sumout ),
	.cout(Xd_0__inst_inst_add_0_98 ),
	.shareout(Xd_0__inst_inst_add_0_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_101 (
// Equation(s):
// Xd_0__inst_inst_add_2_101_sumout  = SUM(( !Xd_0__inst_r_sum1_5__23__q  $ (!Xd_0__inst_r_sum1_4__23__q  $ (Xd_0__inst_r_sum1_3__23__q )) ) + ( Xd_0__inst_inst_add_2_99  ) + ( Xd_0__inst_inst_add_2_98  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__23__q ),
	.datac(!Xd_0__inst_r_sum1_4__23__q ),
	.datad(!Xd_0__inst_r_sum1_3__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_98 ),
	.sharein(Xd_0__inst_inst_add_2_99 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_101_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_101 (
// Equation(s):
// Xd_0__inst_inst_add_0_101_sumout  = SUM(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_99  ) + ( Xd_0__inst_inst_add_0_98  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__23__q ),
	.datad(!Xd_0__inst_r_sum1_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_98 ),
	.sharein(Xd_0__inst_inst_add_0_99 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_101_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_172 (
// Equation(s):
// Xd_0__inst_mult_14_173  = SUM(( GND ) + ( Xd_0__inst_mult_14_179  ) + ( Xd_0__inst_mult_14_178  ))
// Xd_0__inst_mult_14_174  = CARRY(( GND ) + ( Xd_0__inst_mult_14_179  ) + ( Xd_0__inst_mult_14_178  ))
// Xd_0__inst_mult_14_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_178 ),
	.sharein(Xd_0__inst_mult_14_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_173 ),
	.cout(Xd_0__inst_mult_14_174 ),
	.shareout(Xd_0__inst_mult_14_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_172 (
// Equation(s):
// Xd_0__inst_mult_15_173  = SUM(( GND ) + ( Xd_0__inst_mult_15_179  ) + ( Xd_0__inst_mult_15_178  ))
// Xd_0__inst_mult_15_174  = CARRY(( GND ) + ( Xd_0__inst_mult_15_179  ) + ( Xd_0__inst_mult_15_178  ))
// Xd_0__inst_mult_15_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_178 ),
	.sharein(Xd_0__inst_mult_15_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_173 ),
	.cout(Xd_0__inst_mult_15_174 ),
	.shareout(Xd_0__inst_mult_15_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_168 (
// Equation(s):
// Xd_0__inst_mult_12_169  = SUM(( GND ) + ( Xd_0__inst_mult_12_175  ) + ( Xd_0__inst_mult_12_174  ))
// Xd_0__inst_mult_12_170  = CARRY(( GND ) + ( Xd_0__inst_mult_12_175  ) + ( Xd_0__inst_mult_12_174  ))
// Xd_0__inst_mult_12_171  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_174 ),
	.sharein(Xd_0__inst_mult_12_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_169 ),
	.cout(Xd_0__inst_mult_12_170 ),
	.shareout(Xd_0__inst_mult_12_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_70 (
// Equation(s):
// Xd_0__inst_mult_4_180  = SUM(( (!din_a[56] & (((din_a[55] & din_b[58])))) # (din_a[56] & (!din_b[57] $ (((!din_a[55]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_186  ) + ( Xd_0__inst_mult_4_185  ))
// Xd_0__inst_mult_4_181  = CARRY(( (!din_a[56] & (((din_a[55] & din_b[58])))) # (din_a[56] & (!din_b[57] $ (((!din_a[55]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_186  ) + ( Xd_0__inst_mult_4_185  ))
// Xd_0__inst_mult_4_182  = SHARE((din_a[56] & (din_b[57] & (din_a[55] & din_b[58]))))

	.dataa(!din_a[56]),
	.datab(!din_b[57]),
	.datac(!din_a[55]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_185 ),
	.sharein(Xd_0__inst_mult_4_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_180 ),
	.cout(Xd_0__inst_mult_4_181 ),
	.shareout(Xd_0__inst_mult_4_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_12__0__q  $ (!Xd_0__inst_product_13__0__q ) ) + ( Xd_0__inst_mult_9_171  ) + ( Xd_0__inst_mult_9_170  ))
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_12__0__q  $ (!Xd_0__inst_product_13__0__q ) ) + ( Xd_0__inst_mult_9_171  ) + ( Xd_0__inst_mult_9_170  ))
// Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_12__0__q  & ((!Xd_0__inst_sign [13] & ((Xd_0__inst_sign [12]))) # (Xd_0__inst_sign [13] & (!Xd_0__inst_product_13__0__q )))) # (Xd_0__inst_product_12__0__q  & ((!Xd_0__inst_sign [13] 
// & (Xd_0__inst_product_13__0__q )) # (Xd_0__inst_sign [13] & ((!Xd_0__inst_sign [12]))))))

	.dataa(!Xd_0__inst_product_12__0__q ),
	.datab(!Xd_0__inst_product_13__0__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_170 ),
	.sharein(Xd_0__inst_mult_9_171 ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_14__0__q  $ (!Xd_0__inst_product_15__0__q ) ) + ( Xd_0__inst_mult_6_171  ) + ( Xd_0__inst_mult_6_170  ))
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_14__0__q  $ (!Xd_0__inst_product_15__0__q ) ) + ( Xd_0__inst_mult_6_171  ) + ( Xd_0__inst_mult_6_170  ))
// Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_14__0__q  & ((!Xd_0__inst_sign [15] & ((Xd_0__inst_sign [14]))) # (Xd_0__inst_sign [15] & (!Xd_0__inst_product_15__0__q )))) # (Xd_0__inst_product_14__0__q  & ((!Xd_0__inst_sign [15] 
// & (Xd_0__inst_product_15__0__q )) # (Xd_0__inst_sign [15] & ((!Xd_0__inst_sign [14]))))))

	.dataa(!Xd_0__inst_product_14__0__q ),
	.datab(!Xd_0__inst_product_15__0__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_170 ),
	.sharein(Xd_0__inst_mult_6_171 ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14 (
// Equation(s):
// Xd_0__inst_mult_14_177  = SUM(( !Xd_0__inst_mult_14_180  $ (((!din_b[172]) # (!din_a[178]))) ) + ( Xd_0__inst_mult_14_186  ) + ( Xd_0__inst_mult_14_185  ))
// Xd_0__inst_mult_14_178  = CARRY(( !Xd_0__inst_mult_14_180  $ (((!din_b[172]) # (!din_a[178]))) ) + ( Xd_0__inst_mult_14_186  ) + ( Xd_0__inst_mult_14_185  ))
// Xd_0__inst_mult_14_179  = SHARE((din_b[172] & (din_a[178] & Xd_0__inst_mult_14_180 )))

	.dataa(!din_b[172]),
	.datab(!din_a[178]),
	.datac(!Xd_0__inst_mult_14_180 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_185 ),
	.sharein(Xd_0__inst_mult_14_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_177 ),
	.cout(Xd_0__inst_mult_14_178 ),
	.shareout(Xd_0__inst_mult_14_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_10__0__q  $ (!Xd_0__inst_product_11__0__q ) ) + ( Xd_0__inst_mult_8_175  ) + ( Xd_0__inst_mult_8_174  ))
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_10__0__q  $ (!Xd_0__inst_product_11__0__q ) ) + ( Xd_0__inst_mult_8_175  ) + ( Xd_0__inst_mult_8_174  ))
// Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_10__0__q  & ((!Xd_0__inst_sign [11] & ((Xd_0__inst_sign [10]))) # (Xd_0__inst_sign [11] & (!Xd_0__inst_product_11__0__q )))) # (Xd_0__inst_product_10__0__q  & ((!Xd_0__inst_sign [11] 
// & (Xd_0__inst_product_11__0__q )) # (Xd_0__inst_sign [11] & ((!Xd_0__inst_sign [10]))))))

	.dataa(!Xd_0__inst_product_10__0__q ),
	.datab(!Xd_0__inst_product_11__0__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_174 ),
	.sharein(Xd_0__inst_mult_8_175 ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_8__0__q  $ (!Xd_0__inst_product_9__0__q ) ) + ( Xd_0__inst_mult_11_175  ) + ( Xd_0__inst_mult_11_174  ))
// Xd_0__inst_a1_4__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_8__0__q  $ (!Xd_0__inst_product_9__0__q ) ) + ( Xd_0__inst_mult_11_175  ) + ( Xd_0__inst_mult_11_174  ))
// Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_8__0__q  & ((!Xd_0__inst_sign [9] & ((Xd_0__inst_sign [8]))) # (Xd_0__inst_sign [9] & (!Xd_0__inst_product_9__0__q )))) # (Xd_0__inst_product_8__0__q  & ((!Xd_0__inst_sign [9] & 
// (Xd_0__inst_product_9__0__q )) # (Xd_0__inst_sign [9] & ((!Xd_0__inst_sign [8]))))))

	.dataa(!Xd_0__inst_product_8__0__q ),
	.datab(!Xd_0__inst_product_9__0__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_174 ),
	.sharein(Xd_0__inst_mult_11_175 ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( Xd_0__inst_mult_10_171  ) + ( Xd_0__inst_mult_10_170  ))
// Xd_0__inst_a1_3__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( Xd_0__inst_mult_10_171  ) + ( Xd_0__inst_mult_10_170  ))
// Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & ((Xd_0__inst_sign [6]))) # (Xd_0__inst_sign [7] & (!Xd_0__inst_product_7__0__q )))) # (Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & 
// (Xd_0__inst_product_7__0__q )) # (Xd_0__inst_sign [7] & ((!Xd_0__inst_sign [6]))))))

	.dataa(!Xd_0__inst_product_6__0__q ),
	.datab(!Xd_0__inst_product_7__0__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_170 ),
	.sharein(Xd_0__inst_mult_10_171 ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15 (
// Equation(s):
// Xd_0__inst_mult_15_177  = SUM(( (din_a[188] & din_b[190]) ) + ( Xd_0__inst_mult_15_182  ) + ( Xd_0__inst_mult_15_181  ))
// Xd_0__inst_mult_15_178  = CARRY(( (din_a[188] & din_b[190]) ) + ( Xd_0__inst_mult_15_182  ) + ( Xd_0__inst_mult_15_181  ))
// Xd_0__inst_mult_15_179  = SHARE(GND)

	.dataa(!din_a[188]),
	.datab(!din_b[190]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_181 ),
	.sharein(Xd_0__inst_mult_15_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_177 ),
	.cout(Xd_0__inst_mult_15_178 ),
	.shareout(Xd_0__inst_mult_15_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( Xd_0__inst_mult_13_175  ) + ( Xd_0__inst_mult_13_174  ))
// Xd_0__inst_a1_2__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( Xd_0__inst_mult_13_175  ) + ( Xd_0__inst_mult_13_174  ))
// Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & ((Xd_0__inst_sign [4]))) # (Xd_0__inst_sign [5] & (!Xd_0__inst_product_5__0__q )))) # (Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & 
// (Xd_0__inst_product_5__0__q )) # (Xd_0__inst_sign [5] & ((!Xd_0__inst_sign [4]))))))

	.dataa(!Xd_0__inst_product_4__0__q ),
	.datab(!Xd_0__inst_product_5__0__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_174 ),
	.sharein(Xd_0__inst_mult_13_175 ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( Xd_0__inst_mult_15_186  ) + ( Xd_0__inst_mult_15_185  ))
// Xd_0__inst_a1_1__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( Xd_0__inst_mult_15_186  ) + ( Xd_0__inst_mult_15_185  ))
// Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & ((Xd_0__inst_sign [2]))) # (Xd_0__inst_sign [3] & (!Xd_0__inst_product_3__0__q )))) # (Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & 
// (Xd_0__inst_product_3__0__q )) # (Xd_0__inst_sign [3] & ((!Xd_0__inst_sign [2]))))))

	.dataa(!Xd_0__inst_product_2__0__q ),
	.datab(!Xd_0__inst_product_3__0__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_185 ),
	.sharein(Xd_0__inst_mult_15_186 ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( Xd_0__inst_mult_12_178  ) + ( Xd_0__inst_mult_12_177  ))
// Xd_0__inst_a1_0__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( Xd_0__inst_mult_12_178  ) + ( Xd_0__inst_mult_12_177  ))
// Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & ((Xd_0__inst_sign [0]))) # (Xd_0__inst_sign [1] & (!Xd_0__inst_product_1__0__q )))) # (Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & 
// (Xd_0__inst_product_1__0__q )) # (Xd_0__inst_sign [1] & ((!Xd_0__inst_sign [0]))))))

	.dataa(!Xd_0__inst_product_0__0__q ),
	.datab(!Xd_0__inst_product_1__0__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_177 ),
	.sharein(Xd_0__inst_mult_12_178 ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12 (
// Equation(s):
// Xd_0__inst_mult_12_173  = SUM(( (din_a[152] & din_b[154]) ) + ( Xd_0__inst_mult_12_182  ) + ( Xd_0__inst_mult_12_181  ))
// Xd_0__inst_mult_12_174  = CARRY(( (din_a[152] & din_b[154]) ) + ( Xd_0__inst_mult_12_182  ) + ( Xd_0__inst_mult_12_181  ))
// Xd_0__inst_mult_12_175  = SHARE(GND)

	.dataa(!din_a[152]),
	.datab(!din_b[154]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_181 ),
	.sharein(Xd_0__inst_mult_12_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_173 ),
	.cout(Xd_0__inst_mult_12_174 ),
	.shareout(Xd_0__inst_mult_12_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_71 (
// Equation(s):
// Xd_0__inst_mult_4_184  = SUM(( (!din_a[55] & (((din_a[54] & din_b[58])))) # (din_a[55] & (!din_b[57] $ (((!din_a[54]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_190  ) + ( Xd_0__inst_mult_4_189  ))
// Xd_0__inst_mult_4_185  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[58])))) # (din_a[55] & (!din_b[57] $ (((!din_a[54]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_190  ) + ( Xd_0__inst_mult_4_189  ))
// Xd_0__inst_mult_4_186  = SHARE((din_a[55] & (din_b[57] & (din_a[54] & din_b[58]))))

	.dataa(!din_a[55]),
	.datab(!din_b[57]),
	.datac(!din_a[54]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_189 ),
	.sharein(Xd_0__inst_mult_4_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_184 ),
	.cout(Xd_0__inst_mult_4_185 ),
	.shareout(Xd_0__inst_mult_4_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_12__1__q  $ (!Xd_0__inst_product_13__1__q  $ (((Xd_0__inst_sign [13]) # (Xd_0__inst_sign [12])))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_12__1__q  $ (!Xd_0__inst_product_13__1__q  $ (((Xd_0__inst_sign [13]) # (Xd_0__inst_sign [12])))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [12] & (Xd_0__inst_product_12__1__q  & (!Xd_0__inst_product_13__1__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_sign [12] & ((!Xd_0__inst_product_13__1__q  & ((Xd_0__inst_sign [13]))) # 
// (Xd_0__inst_product_13__1__q  & (!Xd_0__inst_product_12__1__q )))))

	.dataa(!Xd_0__inst_product_12__1__q ),
	.datab(!Xd_0__inst_product_13__1__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_14__1__q  $ (!Xd_0__inst_product_15__1__q  $ (((Xd_0__inst_sign [15]) # (Xd_0__inst_sign [14])))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_14__1__q  $ (!Xd_0__inst_product_15__1__q  $ (((Xd_0__inst_sign [15]) # (Xd_0__inst_sign [14])))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [14] & (Xd_0__inst_product_14__1__q  & (!Xd_0__inst_product_15__1__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_sign [14] & ((!Xd_0__inst_product_15__1__q  & ((Xd_0__inst_sign [15]))) # 
// (Xd_0__inst_product_15__1__q  & (!Xd_0__inst_product_14__1__q )))))

	.dataa(!Xd_0__inst_product_14__1__q ),
	.datab(!Xd_0__inst_product_15__1__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_10__1__q  $ (!Xd_0__inst_product_11__1__q  $ (((Xd_0__inst_sign [11]) # (Xd_0__inst_sign [10])))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_10__1__q  $ (!Xd_0__inst_product_11__1__q  $ (((Xd_0__inst_sign [11]) # (Xd_0__inst_sign [10])))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [10] & (Xd_0__inst_product_10__1__q  & (!Xd_0__inst_product_11__1__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_sign [10] & ((!Xd_0__inst_product_11__1__q  & ((Xd_0__inst_sign [11]))) # 
// (Xd_0__inst_product_11__1__q  & (!Xd_0__inst_product_10__1__q )))))

	.dataa(!Xd_0__inst_product_10__1__q ),
	.datab(!Xd_0__inst_product_11__1__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_8__1__q  $ (!Xd_0__inst_product_9__1__q  $ (((Xd_0__inst_sign [9]) # (Xd_0__inst_sign [8])))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_4__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_8__1__q  $ (!Xd_0__inst_product_9__1__q  $ (((Xd_0__inst_sign [9]) # (Xd_0__inst_sign [8])))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [8] & (Xd_0__inst_product_8__1__q  & (!Xd_0__inst_product_9__1__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_sign [8] & ((!Xd_0__inst_product_9__1__q  & ((Xd_0__inst_sign [9]))) # 
// (Xd_0__inst_product_9__1__q  & (!Xd_0__inst_product_8__1__q )))))

	.dataa(!Xd_0__inst_product_8__1__q ),
	.datab(!Xd_0__inst_product_9__1__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [6] & (Xd_0__inst_product_6__1__q  & (!Xd_0__inst_product_7__1__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_sign [6] & ((!Xd_0__inst_product_7__1__q  & ((Xd_0__inst_sign [7]))) # 
// (Xd_0__inst_product_7__1__q  & (!Xd_0__inst_product_6__1__q )))))

	.dataa(!Xd_0__inst_product_6__1__q ),
	.datab(!Xd_0__inst_product_7__1__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [4] & (Xd_0__inst_product_4__1__q  & (!Xd_0__inst_product_5__1__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_sign [4] & ((!Xd_0__inst_product_5__1__q  & ((Xd_0__inst_sign [5]))) # 
// (Xd_0__inst_product_5__1__q  & (!Xd_0__inst_product_4__1__q )))))

	.dataa(!Xd_0__inst_product_4__1__q ),
	.datab(!Xd_0__inst_product_5__1__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [2] & (Xd_0__inst_product_2__1__q  & (!Xd_0__inst_product_3__1__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_sign [2] & ((!Xd_0__inst_product_3__1__q  & ((Xd_0__inst_sign [3]))) # 
// (Xd_0__inst_product_3__1__q  & (!Xd_0__inst_product_2__1__q )))))

	.dataa(!Xd_0__inst_product_2__1__q ),
	.datab(!Xd_0__inst_product_3__1__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [0] & (Xd_0__inst_product_0__1__q  & (!Xd_0__inst_product_1__1__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_sign [0] & ((!Xd_0__inst_product_1__1__q  & ((Xd_0__inst_sign [1]))) # 
// (Xd_0__inst_product_1__1__q  & (!Xd_0__inst_product_0__1__q )))))

	.dataa(!Xd_0__inst_product_0__1__q ),
	.datab(!Xd_0__inst_product_1__1__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_12__2__q  $ (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_12__2__q  $ (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__2__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__2__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__2__q ),
	.datab(!Xd_0__inst_product_13__2__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_14__2__q  $ (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_14__2__q  $ (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__2__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__2__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__2__q ),
	.datab(!Xd_0__inst_product_15__2__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_10__2__q  $ (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_10__2__q  $ (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__2__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__2__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__2__q ),
	.datab(!Xd_0__inst_product_11__2__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_8__2__q  $ (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_8__2__q  $ (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__2__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__2__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__2__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__2__q ),
	.datab(!Xd_0__inst_product_9__2__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__2__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__2__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__2__q ),
	.datab(!Xd_0__inst_product_7__2__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__2__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__2__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__2__q ),
	.datab(!Xd_0__inst_product_5__2__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__2__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__2__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__2__q ),
	.datab(!Xd_0__inst_product_3__2__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__2__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__2__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__2__q ),
	.datab(!Xd_0__inst_product_1__2__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_12__3__q  $ (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_12__3__q  $ (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__3__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__3__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__3__q ),
	.datab(!Xd_0__inst_product_13__3__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_14__3__q  $ (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_14__3__q  $ (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__3__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__3__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__3__q ),
	.datab(!Xd_0__inst_product_15__3__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_10__3__q  $ (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_10__3__q  $ (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__3__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__3__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__3__q ),
	.datab(!Xd_0__inst_product_11__3__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_8__3__q  $ (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_8__3__q  $ (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__3__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__3__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__3__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__3__q ),
	.datab(!Xd_0__inst_product_9__3__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__3__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__3__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__3__q ),
	.datab(!Xd_0__inst_product_7__3__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__3__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__3__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__3__q ),
	.datab(!Xd_0__inst_product_5__3__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__3__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__3__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__3__q ),
	.datab(!Xd_0__inst_product_3__3__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__3__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__3__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__3__q ),
	.datab(!Xd_0__inst_product_1__3__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_12__4__q  $ (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_12__4__q  $ (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__4__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__4__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__4__q ),
	.datab(!Xd_0__inst_product_13__4__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_14__4__q  $ (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_14__4__q  $ (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__4__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__4__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__4__q ),
	.datab(!Xd_0__inst_product_15__4__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_10__4__q  $ (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_10__4__q  $ (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__4__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__4__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__4__q ),
	.datab(!Xd_0__inst_product_11__4__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_8__4__q  $ (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_8__4__q  $ (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__4__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__4__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__4__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__4__q ),
	.datab(!Xd_0__inst_product_9__4__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__4__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__4__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__4__q ),
	.datab(!Xd_0__inst_product_7__4__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__4__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__4__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__4__q ),
	.datab(!Xd_0__inst_product_5__4__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__4__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__4__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__4__q ),
	.datab(!Xd_0__inst_product_3__4__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__4__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__4__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__4__q ),
	.datab(!Xd_0__inst_product_1__4__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_12__5__q  $ (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_12__5__q  $ (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__5__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__5__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__5__q ),
	.datab(!Xd_0__inst_product_13__5__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_14__5__q  $ (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_14__5__q  $ (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__5__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__5__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__5__q ),
	.datab(!Xd_0__inst_product_15__5__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_10__5__q  $ (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_10__5__q  $ (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__5__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__5__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__5__q ),
	.datab(!Xd_0__inst_product_11__5__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_8__5__q  $ (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_8__5__q  $ (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__5__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__5__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__5__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__5__q ),
	.datab(!Xd_0__inst_product_9__5__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__5__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__5__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__5__q ),
	.datab(!Xd_0__inst_product_7__5__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__5__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__5__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__5__q ),
	.datab(!Xd_0__inst_product_5__5__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__5__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__5__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__5__q ),
	.datab(!Xd_0__inst_product_3__5__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__5__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__5__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__5__q ),
	.datab(!Xd_0__inst_product_1__5__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_12__6__q  $ (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_12__6__q  $ (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__6__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__6__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__6__q ),
	.datab(!Xd_0__inst_product_13__6__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_14__6__q  $ (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_14__6__q  $ (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__6__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__6__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__6__q ),
	.datab(!Xd_0__inst_product_15__6__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_10__6__q  $ (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_10__6__q  $ (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__6__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__6__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__6__q ),
	.datab(!Xd_0__inst_product_11__6__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_8__6__q  $ (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_8__6__q  $ (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__6__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__6__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__6__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__6__q ),
	.datab(!Xd_0__inst_product_9__6__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__6__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__6__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__6__q ),
	.datab(!Xd_0__inst_product_7__6__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__6__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__6__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__6__q ),
	.datab(!Xd_0__inst_product_5__6__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__6__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__6__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__6__q ),
	.datab(!Xd_0__inst_product_3__6__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__6__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__6__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__6__q ),
	.datab(!Xd_0__inst_product_1__6__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_12__7__q  $ (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_12__7__q  $ (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__7__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__7__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__7__q ),
	.datab(!Xd_0__inst_product_13__7__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_14__7__q  $ (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_14__7__q  $ (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__7__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__7__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__7__q ),
	.datab(!Xd_0__inst_product_15__7__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_10__7__q  $ (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_10__7__q  $ (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__7__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__7__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__7__q ),
	.datab(!Xd_0__inst_product_11__7__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_8__7__q  $ (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_8__7__q  $ (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__7__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__7__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__7__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__7__q ),
	.datab(!Xd_0__inst_product_9__7__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__7__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__7__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__7__q ),
	.datab(!Xd_0__inst_product_7__7__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__7__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__7__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__7__q ),
	.datab(!Xd_0__inst_product_5__7__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__7__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__7__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__7__q ),
	.datab(!Xd_0__inst_product_3__7__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__7__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__7__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__7__q ),
	.datab(!Xd_0__inst_product_1__7__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_12__8__q  $ (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_12__8__q  $ (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__8__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__8__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__8__q ),
	.datab(!Xd_0__inst_product_13__8__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_14__8__q  $ (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_14__8__q  $ (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__8__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__8__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__8__q ),
	.datab(!Xd_0__inst_product_15__8__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_10__8__q  $ (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_10__8__q  $ (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__8__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__8__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__8__q ),
	.datab(!Xd_0__inst_product_11__8__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_8__8__q  $ (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_8__8__q  $ (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__8__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__8__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__8__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__8__q ),
	.datab(!Xd_0__inst_product_9__8__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__8__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__8__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__8__q ),
	.datab(!Xd_0__inst_product_7__8__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__8__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__8__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__8__q ),
	.datab(!Xd_0__inst_product_5__8__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__8__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__8__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__8__q ),
	.datab(!Xd_0__inst_product_3__8__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__8__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__8__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__8__q ),
	.datab(!Xd_0__inst_product_1__8__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_12__9__q  $ (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_12__9__q  $ (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__9__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__9__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__9__q ),
	.datab(!Xd_0__inst_product_13__9__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_14__9__q  $ (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_14__9__q  $ (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__9__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__9__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__9__q ),
	.datab(!Xd_0__inst_product_15__9__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_10__9__q  $ (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_10__9__q  $ (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__9__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__9__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__9__q ),
	.datab(!Xd_0__inst_product_11__9__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_8__9__q  $ (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_8__9__q  $ (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__9__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__9__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__9__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__9__q ),
	.datab(!Xd_0__inst_product_9__9__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__9__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__9__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__9__q ),
	.datab(!Xd_0__inst_product_7__9__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__9__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__9__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__9__q ),
	.datab(!Xd_0__inst_product_5__9__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__9__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__9__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__9__q ),
	.datab(!Xd_0__inst_product_3__9__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__9__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__9__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__9__q ),
	.datab(!Xd_0__inst_product_1__9__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_12__10__q  $ (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_12__10__q  $ (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__10__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__10__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__10__q ),
	.datab(!Xd_0__inst_product_13__10__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_14__10__q  $ (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_14__10__q  $ (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__10__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__10__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__10__q ),
	.datab(!Xd_0__inst_product_15__10__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_10__10__q  $ (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_10__10__q  $ (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__10__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__10__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__10__q ),
	.datab(!Xd_0__inst_product_11__10__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_8__10__q  $ (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_8__10__q  $ (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__10__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__10__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__10__q ),
	.datab(!Xd_0__inst_product_9__10__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_6__10__q  $ (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_6__10__q  $ (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__10__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__10__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__10__q ),
	.datab(!Xd_0__inst_product_7__10__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_4__10__q  $ (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_4__10__q  $ (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__10__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__10__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__10__q ),
	.datab(!Xd_0__inst_product_5__10__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_2__10__q  $ (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_2__10__q  $ (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__10__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__10__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__10__q ),
	.datab(!Xd_0__inst_product_3__10__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_0__10__q  $ (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_0__10__q  $ (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__10__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__10__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__10__q ),
	.datab(!Xd_0__inst_product_1__10__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_12__11__q  $ (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_12__11__q  $ (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__11__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__11__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__11__q ),
	.datab(!Xd_0__inst_product_13__11__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_14__11__q  $ (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_14__11__q  $ (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__11__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__11__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__11__q ),
	.datab(!Xd_0__inst_product_15__11__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_10__11__q  $ (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_10__11__q  $ (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__11__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__11__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__11__q ),
	.datab(!Xd_0__inst_product_11__11__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_8__11__q  $ (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_8__11__q  $ (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__11__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__11__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__11__q ),
	.datab(!Xd_0__inst_product_9__11__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_6__11__q  $ (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_6__11__q  $ (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__11__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__11__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__11__q ),
	.datab(!Xd_0__inst_product_7__11__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_4__11__q  $ (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_4__11__q  $ (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__11__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__11__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__11__q ),
	.datab(!Xd_0__inst_product_5__11__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_2__11__q  $ (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_2__11__q  $ (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__11__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__11__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__11__q ),
	.datab(!Xd_0__inst_product_3__11__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_0__11__q  $ (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_0__11__q  $ (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__11__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__11__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__11__q ),
	.datab(!Xd_0__inst_product_1__11__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_12__12__q  $ (!Xd_0__inst_product_13__12__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_12__12__q  $ (!Xd_0__inst_product_13__12__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__12__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__12__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__12__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__12__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__12__q ),
	.datab(!Xd_0__inst_product_13__12__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_14__12__q  $ (!Xd_0__inst_product_15__12__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_14__12__q  $ (!Xd_0__inst_product_15__12__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__12__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__12__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__12__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__12__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__12__q ),
	.datab(!Xd_0__inst_product_15__12__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_10__12__q  $ (!Xd_0__inst_product_11__12__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_10__12__q  $ (!Xd_0__inst_product_11__12__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__12__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__12__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__12__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__12__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__12__q ),
	.datab(!Xd_0__inst_product_11__12__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_8__12__q  $ (!Xd_0__inst_product_9__12__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_8__12__q  $ (!Xd_0__inst_product_9__12__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__12__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__12__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__12__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__12__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__12__q ),
	.datab(!Xd_0__inst_product_9__12__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_6__12__q  $ (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_6__12__q  $ (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__12__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__12__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__12__q ),
	.datab(!Xd_0__inst_product_7__12__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_4__12__q  $ (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_4__12__q  $ (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__12__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__12__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__12__q ),
	.datab(!Xd_0__inst_product_5__12__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_2__12__q  $ (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_2__12__q  $ (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__12__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__12__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__12__q ),
	.datab(!Xd_0__inst_product_3__12__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_0__12__q  $ (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_0__12__q  $ (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__12__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__12__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__12__q ),
	.datab(!Xd_0__inst_product_1__12__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_12__13__q  $ (!Xd_0__inst_product_13__13__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_12__13__q  $ (!Xd_0__inst_product_13__13__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__13__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__13__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__13__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__13__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__13__q ),
	.datab(!Xd_0__inst_product_13__13__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_14__13__q  $ (!Xd_0__inst_product_15__13__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_14__13__q  $ (!Xd_0__inst_product_15__13__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__13__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__13__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__13__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__13__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__13__q ),
	.datab(!Xd_0__inst_product_15__13__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_10__13__q  $ (!Xd_0__inst_product_11__13__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_10__13__q  $ (!Xd_0__inst_product_11__13__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__13__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__13__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__13__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__13__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__13__q ),
	.datab(!Xd_0__inst_product_11__13__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_8__13__q  $ (!Xd_0__inst_product_9__13__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_8__13__q  $ (!Xd_0__inst_product_9__13__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__13__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__13__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__13__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__13__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__13__q ),
	.datab(!Xd_0__inst_product_9__13__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_6__13__q  $ (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_6__13__q  $ (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__13__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__13__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__13__q ),
	.datab(!Xd_0__inst_product_7__13__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_4__13__q  $ (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_4__13__q  $ (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__13__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__13__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__13__q ),
	.datab(!Xd_0__inst_product_5__13__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_2__13__q  $ (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_2__13__q  $ (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__13__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__13__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__13__q ),
	.datab(!Xd_0__inst_product_3__13__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_0__13__q  $ (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_0__13__q  $ (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__13__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__13__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__13__q ),
	.datab(!Xd_0__inst_product_1__13__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_12__14__q  $ (!Xd_0__inst_product_13__14__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_12__14__q  $ (!Xd_0__inst_product_13__14__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__14__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__14__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__14__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__14__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__14__q ),
	.datab(!Xd_0__inst_product_13__14__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_14__14__q  $ (!Xd_0__inst_product_15__14__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_14__14__q  $ (!Xd_0__inst_product_15__14__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__14__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__14__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__14__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__14__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__14__q ),
	.datab(!Xd_0__inst_product_15__14__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_10__14__q  $ (!Xd_0__inst_product_11__14__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_10__14__q  $ (!Xd_0__inst_product_11__14__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__14__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__14__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__14__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__14__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__14__q ),
	.datab(!Xd_0__inst_product_11__14__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_8__14__q  $ (!Xd_0__inst_product_9__14__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_8__14__q  $ (!Xd_0__inst_product_9__14__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__14__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__14__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__14__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__14__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__14__q ),
	.datab(!Xd_0__inst_product_9__14__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_6__14__q  $ (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_6__14__q  $ (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__14__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__14__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__14__q ),
	.datab(!Xd_0__inst_product_7__14__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_4__14__q  $ (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_4__14__q  $ (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__14__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__14__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__14__q ),
	.datab(!Xd_0__inst_product_5__14__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_2__14__q  $ (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_2__14__q  $ (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__14__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__14__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__14__q ),
	.datab(!Xd_0__inst_product_3__14__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_0__14__q  $ (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_0__14__q  $ (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__14__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__14__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__14__q ),
	.datab(!Xd_0__inst_product_1__14__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_12__15__q  $ (!Xd_0__inst_product_13__15__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_12__15__q  $ (!Xd_0__inst_product_13__15__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__15__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__15__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__15__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__15__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__15__q ),
	.datab(!Xd_0__inst_product_13__15__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_14__15__q  $ (!Xd_0__inst_product_15__15__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_14__15__q  $ (!Xd_0__inst_product_15__15__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__15__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__15__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__15__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__15__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__15__q ),
	.datab(!Xd_0__inst_product_15__15__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_10__15__q  $ (!Xd_0__inst_product_11__15__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_10__15__q  $ (!Xd_0__inst_product_11__15__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__15__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__15__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__15__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__15__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__15__q ),
	.datab(!Xd_0__inst_product_11__15__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_8__15__q  $ (!Xd_0__inst_product_9__15__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_8__15__q  $ (!Xd_0__inst_product_9__15__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__15__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__15__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__15__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__15__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__15__q ),
	.datab(!Xd_0__inst_product_9__15__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_6__15__q  $ (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_6__15__q  $ (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__15__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__15__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__15__q ),
	.datab(!Xd_0__inst_product_7__15__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_4__15__q  $ (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_4__15__q  $ (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__15__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__15__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__15__q ),
	.datab(!Xd_0__inst_product_5__15__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_2__15__q  $ (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_2__15__q  $ (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__15__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__15__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__15__q ),
	.datab(!Xd_0__inst_product_3__15__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_0__15__q  $ (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_0__15__q  $ (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__15__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__15__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__15__q ),
	.datab(!Xd_0__inst_product_1__15__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_12__16__q  $ (!Xd_0__inst_product_13__16__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_12__16__q  $ (!Xd_0__inst_product_13__16__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__16__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__16__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__16__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__16__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__16__q ),
	.datab(!Xd_0__inst_product_13__16__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_14__16__q  $ (!Xd_0__inst_product_15__16__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_14__16__q  $ (!Xd_0__inst_product_15__16__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__16__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__16__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__16__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__16__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__16__q ),
	.datab(!Xd_0__inst_product_15__16__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_10__16__q  $ (!Xd_0__inst_product_11__16__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_10__16__q  $ (!Xd_0__inst_product_11__16__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__16__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__16__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__16__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__16__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__16__q ),
	.datab(!Xd_0__inst_product_11__16__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_8__16__q  $ (!Xd_0__inst_product_9__16__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_8__16__q  $ (!Xd_0__inst_product_9__16__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__16__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__16__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__16__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__16__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__16__q ),
	.datab(!Xd_0__inst_product_9__16__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_6__16__q  $ (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_6__16__q  $ (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__16__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__16__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__16__q ),
	.datab(!Xd_0__inst_product_7__16__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_4__16__q  $ (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_4__16__q  $ (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__16__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__16__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__16__q ),
	.datab(!Xd_0__inst_product_5__16__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_2__16__q  $ (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_2__16__q  $ (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__16__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__16__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__16__q ),
	.datab(!Xd_0__inst_product_3__16__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_0__16__q  $ (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_0__16__q  $ (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__16__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__16__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__16__q ),
	.datab(!Xd_0__inst_product_1__16__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_12__17__q  $ (!Xd_0__inst_product_13__17__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_12__17__q  $ (!Xd_0__inst_product_13__17__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__17__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__17__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__17__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__17__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__17__q ),
	.datab(!Xd_0__inst_product_13__17__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_14__17__q  $ (!Xd_0__inst_product_15__17__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_14__17__q  $ (!Xd_0__inst_product_15__17__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__17__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__17__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__17__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__17__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__17__q ),
	.datab(!Xd_0__inst_product_15__17__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_10__17__q  $ (!Xd_0__inst_product_11__17__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_10__17__q  $ (!Xd_0__inst_product_11__17__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__17__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__17__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__17__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__17__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__17__q ),
	.datab(!Xd_0__inst_product_11__17__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_8__17__q  $ (!Xd_0__inst_product_9__17__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_8__17__q  $ (!Xd_0__inst_product_9__17__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__17__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__17__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__17__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__17__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__17__q ),
	.datab(!Xd_0__inst_product_9__17__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_6__17__q  $ (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_6__17__q  $ (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__17__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__17__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__17__q ),
	.datab(!Xd_0__inst_product_7__17__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_4__17__q  $ (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_4__17__q  $ (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__17__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__17__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__17__q ),
	.datab(!Xd_0__inst_product_5__17__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_2__17__q  $ (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_2__17__q  $ (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__17__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__17__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__17__q ),
	.datab(!Xd_0__inst_product_3__17__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_0__17__q  $ (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_0__17__q  $ (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__17__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__17__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__17__q ),
	.datab(!Xd_0__inst_product_1__17__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_12__18__q  $ (!Xd_0__inst_product_13__18__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_12__18__q  $ (!Xd_0__inst_product_13__18__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__18__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__18__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__18__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__18__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__18__q ),
	.datab(!Xd_0__inst_product_13__18__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_14__18__q  $ (!Xd_0__inst_product_15__18__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_14__18__q  $ (!Xd_0__inst_product_15__18__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__18__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__18__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__18__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__18__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__18__q ),
	.datab(!Xd_0__inst_product_15__18__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_10__18__q  $ (!Xd_0__inst_product_11__18__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_10__18__q  $ (!Xd_0__inst_product_11__18__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__18__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__18__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__18__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__18__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__18__q ),
	.datab(!Xd_0__inst_product_11__18__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_8__18__q  $ (!Xd_0__inst_product_9__18__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_8__18__q  $ (!Xd_0__inst_product_9__18__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__18__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__18__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__18__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__18__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__18__q ),
	.datab(!Xd_0__inst_product_9__18__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_6__18__q  $ (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_6__18__q  $ (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__18__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__18__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__18__q ),
	.datab(!Xd_0__inst_product_7__18__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_4__18__q  $ (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_4__18__q  $ (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__18__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__18__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__18__q ),
	.datab(!Xd_0__inst_product_5__18__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_2__18__q  $ (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_2__18__q  $ (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__18__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__18__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__18__q ),
	.datab(!Xd_0__inst_product_3__18__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_0__18__q  $ (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_0__18__q  $ (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__18__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__18__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__18__q ),
	.datab(!Xd_0__inst_product_1__18__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_12__19__q  $ (!Xd_0__inst_product_13__19__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_12__19__q  $ (!Xd_0__inst_product_13__19__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__19__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__19__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__19__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__19__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__19__q ),
	.datab(!Xd_0__inst_product_13__19__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_14__19__q  $ (!Xd_0__inst_product_15__19__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_14__19__q  $ (!Xd_0__inst_product_15__19__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__19__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__19__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__19__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__19__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__19__q ),
	.datab(!Xd_0__inst_product_15__19__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_10__19__q  $ (!Xd_0__inst_product_11__19__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_10__19__q  $ (!Xd_0__inst_product_11__19__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__19__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__19__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__19__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__19__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__19__q ),
	.datab(!Xd_0__inst_product_11__19__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_8__19__q  $ (!Xd_0__inst_product_9__19__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_8__19__q  $ (!Xd_0__inst_product_9__19__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__19__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__19__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__19__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__19__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__19__q ),
	.datab(!Xd_0__inst_product_9__19__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_6__19__q  $ (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_6__19__q  $ (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__19__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__19__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__19__q ),
	.datab(!Xd_0__inst_product_7__19__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_4__19__q  $ (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_4__19__q  $ (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__19__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__19__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__19__q ),
	.datab(!Xd_0__inst_product_5__19__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_2__19__q  $ (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_2__19__q  $ (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__19__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__19__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__19__q ),
	.datab(!Xd_0__inst_product_3__19__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_0__19__q  $ (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_0__19__q  $ (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__19__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__19__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__19__q ),
	.datab(!Xd_0__inst_product_1__19__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_12__20__q  $ (!Xd_0__inst_product_13__20__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_12__20__q  $ (!Xd_0__inst_product_13__20__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__20__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__20__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__20__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__20__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__20__q ),
	.datab(!Xd_0__inst_product_13__20__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_14__20__q  $ (!Xd_0__inst_product_15__20__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_14__20__q  $ (!Xd_0__inst_product_15__20__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__20__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__20__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__20__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__20__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__20__q ),
	.datab(!Xd_0__inst_product_15__20__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_10__20__q  $ (!Xd_0__inst_product_11__20__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_10__20__q  $ (!Xd_0__inst_product_11__20__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__20__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__20__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__20__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__20__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__20__q ),
	.datab(!Xd_0__inst_product_11__20__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_8__20__q  $ (!Xd_0__inst_product_9__20__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_8__20__q  $ (!Xd_0__inst_product_9__20__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__20__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__20__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__20__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__20__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__20__q ),
	.datab(!Xd_0__inst_product_9__20__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_6__20__q  $ (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_6__20__q  $ (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__20__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__20__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__20__q ),
	.datab(!Xd_0__inst_product_7__20__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_4__20__q  $ (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_4__20__q  $ (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__20__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__20__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__20__q ),
	.datab(!Xd_0__inst_product_5__20__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_2__20__q  $ (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_2__20__q  $ (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__20__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__20__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__20__q ),
	.datab(!Xd_0__inst_product_3__20__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_0__20__q  $ (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_0__20__q  $ (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__20__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__20__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__20__q ),
	.datab(!Xd_0__inst_product_1__20__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_12__21__q  $ (!Xd_0__inst_product_13__21__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_12__21__q  $ (!Xd_0__inst_product_13__21__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__21__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__21__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__21__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__21__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__21__q ),
	.datab(!Xd_0__inst_product_13__21__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_14__21__q  $ (!Xd_0__inst_product_15__21__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_14__21__q  $ (!Xd_0__inst_product_15__21__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__21__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__21__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__21__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__21__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__21__q ),
	.datab(!Xd_0__inst_product_15__21__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_10__21__q  $ (!Xd_0__inst_product_11__21__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_10__21__q  $ (!Xd_0__inst_product_11__21__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__21__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__21__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__21__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__21__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__21__q ),
	.datab(!Xd_0__inst_product_11__21__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_8__21__q  $ (!Xd_0__inst_product_9__21__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_8__21__q  $ (!Xd_0__inst_product_9__21__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__21__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__21__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__21__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__21__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__21__q ),
	.datab(!Xd_0__inst_product_9__21__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_6__21__q  $ (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_6__21__q  $ (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__21__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__21__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__21__q ),
	.datab(!Xd_0__inst_product_7__21__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_4__21__q  $ (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_4__21__q  $ (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__21__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__21__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__21__q ),
	.datab(!Xd_0__inst_product_5__21__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_2__21__q  $ (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_2__21__q  $ (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__21__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__21__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__21__q ),
	.datab(!Xd_0__inst_product_3__21__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_0__21__q  $ (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_0__21__q  $ (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__21__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__21__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__21__q ),
	.datab(!Xd_0__inst_product_1__21__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [12] & Xd_0__inst_sign [13]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [14] & Xd_0__inst_sign [15]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [10] & Xd_0__inst_sign [11]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [8] & Xd_0__inst_sign [9]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [6] & Xd_0__inst_sign [7]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [4] & Xd_0__inst_sign [5]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [2] & Xd_0__inst_sign [3]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [0] & Xd_0__inst_sign [1]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_168 (
// Equation(s):
// Xd_0__inst_mult_9_169  = SUM(( GND ) + ( Xd_0__inst_mult_9_175  ) + ( Xd_0__inst_mult_9_174  ))
// Xd_0__inst_mult_9_170  = CARRY(( GND ) + ( Xd_0__inst_mult_9_175  ) + ( Xd_0__inst_mult_9_174  ))
// Xd_0__inst_mult_9_171  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_174 ),
	.sharein(Xd_0__inst_mult_9_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_169 ),
	.cout(Xd_0__inst_mult_9_170 ),
	.shareout(Xd_0__inst_mult_9_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_168 (
// Equation(s):
// Xd_0__inst_mult_6_169  = SUM(( GND ) + ( Xd_0__inst_mult_6_175  ) + ( Xd_0__inst_mult_6_174  ))
// Xd_0__inst_mult_6_170  = CARRY(( GND ) + ( Xd_0__inst_mult_6_175  ) + ( Xd_0__inst_mult_6_174  ))
// Xd_0__inst_mult_6_171  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_174 ),
	.sharein(Xd_0__inst_mult_6_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_169 ),
	.cout(Xd_0__inst_mult_6_170 ),
	.shareout(Xd_0__inst_mult_6_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_70 (
// Equation(s):
// Xd_0__inst_mult_14_180  = SUM(( GND ) + ( Xd_0__inst_mult_14_190  ) + ( Xd_0__inst_mult_14_189  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_189 ),
	.sharein(Xd_0__inst_mult_14_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_180 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_71 (
// Equation(s):
// Xd_0__inst_mult_14_184  = SUM(( !Xd_0__inst_mult_14_188  $ (((!din_b[171]) # (!din_a[178]))) ) + ( Xd_0__inst_mult_14_194  ) + ( Xd_0__inst_mult_14_193  ))
// Xd_0__inst_mult_14_185  = CARRY(( !Xd_0__inst_mult_14_188  $ (((!din_b[171]) # (!din_a[178]))) ) + ( Xd_0__inst_mult_14_194  ) + ( Xd_0__inst_mult_14_193  ))
// Xd_0__inst_mult_14_186  = SHARE((din_b[171] & (din_a[178] & Xd_0__inst_mult_14_188 )))

	.dataa(!din_b[171]),
	.datab(!din_a[178]),
	.datac(!Xd_0__inst_mult_14_188 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_193 ),
	.sharein(Xd_0__inst_mult_14_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_184 ),
	.cout(Xd_0__inst_mult_14_185 ),
	.shareout(Xd_0__inst_mult_14_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_172 (
// Equation(s):
// Xd_0__inst_mult_8_173  = SUM(( GND ) + ( Xd_0__inst_mult_8_179  ) + ( Xd_0__inst_mult_8_178  ))
// Xd_0__inst_mult_8_174  = CARRY(( GND ) + ( Xd_0__inst_mult_8_179  ) + ( Xd_0__inst_mult_8_178  ))
// Xd_0__inst_mult_8_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_178 ),
	.sharein(Xd_0__inst_mult_8_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_173 ),
	.cout(Xd_0__inst_mult_8_174 ),
	.shareout(Xd_0__inst_mult_8_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_172 (
// Equation(s):
// Xd_0__inst_mult_11_173  = SUM(( GND ) + ( Xd_0__inst_mult_11_179  ) + ( Xd_0__inst_mult_11_178  ))
// Xd_0__inst_mult_11_174  = CARRY(( GND ) + ( Xd_0__inst_mult_11_179  ) + ( Xd_0__inst_mult_11_178  ))
// Xd_0__inst_mult_11_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_178 ),
	.sharein(Xd_0__inst_mult_11_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_173 ),
	.cout(Xd_0__inst_mult_11_174 ),
	.shareout(Xd_0__inst_mult_11_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_168 (
// Equation(s):
// Xd_0__inst_mult_10_169  = SUM(( GND ) + ( Xd_0__inst_mult_10_175  ) + ( Xd_0__inst_mult_10_174  ))
// Xd_0__inst_mult_10_170  = CARRY(( GND ) + ( Xd_0__inst_mult_10_175  ) + ( Xd_0__inst_mult_10_174  ))
// Xd_0__inst_mult_10_171  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_174 ),
	.sharein(Xd_0__inst_mult_10_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_169 ),
	.cout(Xd_0__inst_mult_10_170 ),
	.shareout(Xd_0__inst_mult_10_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_70 (
// Equation(s):
// Xd_0__inst_mult_15_180  = SUM(( (!din_a[188] & (((din_a[187] & din_b[190])))) # (din_a[188] & (!din_b[189] $ (((!din_a[187]) # (!din_b[190]))))) ) + ( Xd_0__inst_mult_15_190  ) + ( Xd_0__inst_mult_15_189  ))
// Xd_0__inst_mult_15_181  = CARRY(( (!din_a[188] & (((din_a[187] & din_b[190])))) # (din_a[188] & (!din_b[189] $ (((!din_a[187]) # (!din_b[190]))))) ) + ( Xd_0__inst_mult_15_190  ) + ( Xd_0__inst_mult_15_189  ))
// Xd_0__inst_mult_15_182  = SHARE((din_a[188] & (din_b[189] & (din_a[187] & din_b[190]))))

	.dataa(!din_a[188]),
	.datab(!din_b[189]),
	.datac(!din_a[187]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_189 ),
	.sharein(Xd_0__inst_mult_15_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_180 ),
	.cout(Xd_0__inst_mult_15_181 ),
	.shareout(Xd_0__inst_mult_15_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_172 (
// Equation(s):
// Xd_0__inst_mult_13_173  = SUM(( GND ) + ( Xd_0__inst_mult_13_179  ) + ( Xd_0__inst_mult_13_178  ))
// Xd_0__inst_mult_13_174  = CARRY(( GND ) + ( Xd_0__inst_mult_13_179  ) + ( Xd_0__inst_mult_13_178  ))
// Xd_0__inst_mult_13_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_178 ),
	.sharein(Xd_0__inst_mult_13_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_173 ),
	.cout(Xd_0__inst_mult_13_174 ),
	.shareout(Xd_0__inst_mult_13_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_71 (
// Equation(s):
// Xd_0__inst_mult_15_184  = SUM(( GND ) + ( Xd_0__inst_mult_15_194  ) + ( Xd_0__inst_mult_15_193  ))
// Xd_0__inst_mult_15_185  = CARRY(( GND ) + ( Xd_0__inst_mult_15_194  ) + ( Xd_0__inst_mult_15_193  ))
// Xd_0__inst_mult_15_186  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_193 ),
	.sharein(Xd_0__inst_mult_15_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_184 ),
	.cout(Xd_0__inst_mult_15_185 ),
	.shareout(Xd_0__inst_mult_15_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_66 (
// Equation(s):
// Xd_0__inst_mult_12_176  = SUM(( GND ) + ( Xd_0__inst_mult_12_186  ) + ( Xd_0__inst_mult_12_185  ))
// Xd_0__inst_mult_12_177  = CARRY(( GND ) + ( Xd_0__inst_mult_12_186  ) + ( Xd_0__inst_mult_12_185  ))
// Xd_0__inst_mult_12_178  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_185 ),
	.sharein(Xd_0__inst_mult_12_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_176 ),
	.cout(Xd_0__inst_mult_12_177 ),
	.shareout(Xd_0__inst_mult_12_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_67 (
// Equation(s):
// Xd_0__inst_mult_12_180  = SUM(( (!din_a[152] & (((din_a[151] & din_b[154])))) # (din_a[152] & (!din_b[153] $ (((!din_a[151]) # (!din_b[154]))))) ) + ( Xd_0__inst_mult_12_190  ) + ( Xd_0__inst_mult_12_189  ))
// Xd_0__inst_mult_12_181  = CARRY(( (!din_a[152] & (((din_a[151] & din_b[154])))) # (din_a[152] & (!din_b[153] $ (((!din_a[151]) # (!din_b[154]))))) ) + ( Xd_0__inst_mult_12_190  ) + ( Xd_0__inst_mult_12_189  ))
// Xd_0__inst_mult_12_182  = SHARE((din_a[152] & (din_b[153] & (din_a[151] & din_b[154]))))

	.dataa(!din_a[152]),
	.datab(!din_b[153]),
	.datac(!din_a[151]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_189 ),
	.sharein(Xd_0__inst_mult_12_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_180 ),
	.cout(Xd_0__inst_mult_12_181 ),
	.shareout(Xd_0__inst_mult_12_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_72 (
// Equation(s):
// Xd_0__inst_mult_4_188  = SUM(( (!din_a[55] & (((din_a[54] & din_b[57])))) # (din_a[55] & (!din_b[56] $ (((!din_a[54]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_4_194  ) + ( Xd_0__inst_mult_4_193  ))
// Xd_0__inst_mult_4_189  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[57])))) # (din_a[55] & (!din_b[56] $ (((!din_a[54]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_4_194  ) + ( Xd_0__inst_mult_4_193  ))
// Xd_0__inst_mult_4_190  = SHARE((din_a[55] & (din_b[56] & (din_a[54] & din_b[57]))))

	.dataa(!din_a[55]),
	.datab(!din_b[56]),
	.datac(!din_a[54]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_193 ),
	.sharein(Xd_0__inst_mult_4_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_188 ),
	.cout(Xd_0__inst_mult_4_189 ),
	.shareout(Xd_0__inst_mult_4_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9 (
// Equation(s):
// Xd_0__inst_mult_9_173  = SUM(( !Xd_0__inst_mult_9_244  $ (((!din_b[112]) # (!din_a[118]))) ) + ( Xd_0__inst_mult_9_250  ) + ( Xd_0__inst_mult_9_249  ))
// Xd_0__inst_mult_9_174  = CARRY(( !Xd_0__inst_mult_9_244  $ (((!din_b[112]) # (!din_a[118]))) ) + ( Xd_0__inst_mult_9_250  ) + ( Xd_0__inst_mult_9_249  ))
// Xd_0__inst_mult_9_175  = SHARE((din_b[112] & (din_a[118] & Xd_0__inst_mult_9_244 )))

	.dataa(!din_b[112]),
	.datab(!din_a[118]),
	.datac(!Xd_0__inst_mult_9_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_249 ),
	.sharein(Xd_0__inst_mult_9_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_173 ),
	.cout(Xd_0__inst_mult_9_174 ),
	.shareout(Xd_0__inst_mult_9_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6 (
// Equation(s):
// Xd_0__inst_mult_6_173  = SUM(( !Xd_0__inst_mult_6_244  $ (((!din_b[76]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_250  ) + ( Xd_0__inst_mult_6_249  ))
// Xd_0__inst_mult_6_174  = CARRY(( !Xd_0__inst_mult_6_244  $ (((!din_b[76]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_250  ) + ( Xd_0__inst_mult_6_249  ))
// Xd_0__inst_mult_6_175  = SHARE((din_b[76] & (din_a[82] & Xd_0__inst_mult_6_244 )))

	.dataa(!din_b[76]),
	.datab(!din_a[82]),
	.datac(!Xd_0__inst_mult_6_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_249 ),
	.sharein(Xd_0__inst_mult_6_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_173 ),
	.cout(Xd_0__inst_mult_6_174 ),
	.shareout(Xd_0__inst_mult_6_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_72 (
// Equation(s):
// Xd_0__inst_mult_14_188  = SUM(( (din_a[177] & din_b[172]) ) + ( Xd_0__inst_mult_14_270  ) + ( Xd_0__inst_mult_14_269  ))
// Xd_0__inst_mult_14_189  = CARRY(( (din_a[177] & din_b[172]) ) + ( Xd_0__inst_mult_14_270  ) + ( Xd_0__inst_mult_14_269  ))
// Xd_0__inst_mult_14_190  = SHARE(GND)

	.dataa(!din_a[177]),
	.datab(!din_b[172]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_269 ),
	.sharein(Xd_0__inst_mult_14_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_188 ),
	.cout(Xd_0__inst_mult_14_189 ),
	.shareout(Xd_0__inst_mult_14_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_73 (
// Equation(s):
// Xd_0__inst_mult_14_192  = SUM(( !Xd_0__inst_mult_14_272  $ (!Xd_0__inst_mult_14_268  $ (((din_b[170] & din_a[178])))) ) + ( Xd_0__inst_mult_14_278  ) + ( Xd_0__inst_mult_14_277  ))
// Xd_0__inst_mult_14_193  = CARRY(( !Xd_0__inst_mult_14_272  $ (!Xd_0__inst_mult_14_268  $ (((din_b[170] & din_a[178])))) ) + ( Xd_0__inst_mult_14_278  ) + ( Xd_0__inst_mult_14_277  ))
// Xd_0__inst_mult_14_194  = SHARE((!Xd_0__inst_mult_14_272  & (Xd_0__inst_mult_14_268  & (din_b[170] & din_a[178]))) # (Xd_0__inst_mult_14_272  & (((din_b[170] & din_a[178])) # (Xd_0__inst_mult_14_268 ))))

	.dataa(!Xd_0__inst_mult_14_272 ),
	.datab(!Xd_0__inst_mult_14_268 ),
	.datac(!din_b[170]),
	.datad(!din_a[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_277 ),
	.sharein(Xd_0__inst_mult_14_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_192 ),
	.cout(Xd_0__inst_mult_14_193 ),
	.shareout(Xd_0__inst_mult_14_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8 (
// Equation(s):
// Xd_0__inst_mult_8_177  = SUM(( !Xd_0__inst_mult_8_248  $ (((!din_b[100]) # (!din_a[106]))) ) + ( Xd_0__inst_mult_8_254  ) + ( Xd_0__inst_mult_8_253  ))
// Xd_0__inst_mult_8_178  = CARRY(( !Xd_0__inst_mult_8_248  $ (((!din_b[100]) # (!din_a[106]))) ) + ( Xd_0__inst_mult_8_254  ) + ( Xd_0__inst_mult_8_253  ))
// Xd_0__inst_mult_8_179  = SHARE((din_b[100] & (din_a[106] & Xd_0__inst_mult_8_248 )))

	.dataa(!din_b[100]),
	.datab(!din_a[106]),
	.datac(!Xd_0__inst_mult_8_248 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_253 ),
	.sharein(Xd_0__inst_mult_8_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_177 ),
	.cout(Xd_0__inst_mult_8_178 ),
	.shareout(Xd_0__inst_mult_8_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11 (
// Equation(s):
// Xd_0__inst_mult_11_177  = SUM(( !Xd_0__inst_mult_11_252  $ (((!din_b[136]) # (!din_a[142]))) ) + ( Xd_0__inst_mult_11_258  ) + ( Xd_0__inst_mult_11_257  ))
// Xd_0__inst_mult_11_178  = CARRY(( !Xd_0__inst_mult_11_252  $ (((!din_b[136]) # (!din_a[142]))) ) + ( Xd_0__inst_mult_11_258  ) + ( Xd_0__inst_mult_11_257  ))
// Xd_0__inst_mult_11_179  = SHARE((din_b[136] & (din_a[142] & Xd_0__inst_mult_11_252 )))

	.dataa(!din_b[136]),
	.datab(!din_a[142]),
	.datac(!Xd_0__inst_mult_11_252 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_257 ),
	.sharein(Xd_0__inst_mult_11_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_177 ),
	.cout(Xd_0__inst_mult_11_178 ),
	.shareout(Xd_0__inst_mult_11_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10 (
// Equation(s):
// Xd_0__inst_mult_10_173  = SUM(( !Xd_0__inst_mult_10_248  $ (((!din_b[124]) # (!din_a[130]))) ) + ( Xd_0__inst_mult_10_254  ) + ( Xd_0__inst_mult_10_253  ))
// Xd_0__inst_mult_10_174  = CARRY(( !Xd_0__inst_mult_10_248  $ (((!din_b[124]) # (!din_a[130]))) ) + ( Xd_0__inst_mult_10_254  ) + ( Xd_0__inst_mult_10_253  ))
// Xd_0__inst_mult_10_175  = SHARE((din_b[124] & (din_a[130] & Xd_0__inst_mult_10_248 )))

	.dataa(!din_b[124]),
	.datab(!din_a[130]),
	.datac(!Xd_0__inst_mult_10_248 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_253 ),
	.sharein(Xd_0__inst_mult_10_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_173 ),
	.cout(Xd_0__inst_mult_10_174 ),
	.shareout(Xd_0__inst_mult_10_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_72 (
// Equation(s):
// Xd_0__inst_mult_15_188  = SUM(( (!din_a[187] & (((din_a[186] & din_b[190])))) # (din_a[187] & (!din_b[189] $ (((!din_a[186]) # (!din_b[190]))))) ) + ( Xd_0__inst_mult_15_270  ) + ( Xd_0__inst_mult_15_269  ))
// Xd_0__inst_mult_15_189  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[190])))) # (din_a[187] & (!din_b[189] $ (((!din_a[186]) # (!din_b[190]))))) ) + ( Xd_0__inst_mult_15_270  ) + ( Xd_0__inst_mult_15_269  ))
// Xd_0__inst_mult_15_190  = SHARE((din_a[187] & (din_b[189] & (din_a[186] & din_b[190]))))

	.dataa(!din_a[187]),
	.datab(!din_b[189]),
	.datac(!din_a[186]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_269 ),
	.sharein(Xd_0__inst_mult_15_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_188 ),
	.cout(Xd_0__inst_mult_15_189 ),
	.shareout(Xd_0__inst_mult_15_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13 (
// Equation(s):
// Xd_0__inst_mult_13_177  = SUM(( !Xd_0__inst_mult_13_252  $ (((!din_b[160]) # (!din_a[166]))) ) + ( Xd_0__inst_mult_13_258  ) + ( Xd_0__inst_mult_13_257  ))
// Xd_0__inst_mult_13_178  = CARRY(( !Xd_0__inst_mult_13_252  $ (((!din_b[160]) # (!din_a[166]))) ) + ( Xd_0__inst_mult_13_258  ) + ( Xd_0__inst_mult_13_257  ))
// Xd_0__inst_mult_13_179  = SHARE((din_b[160] & (din_a[166] & Xd_0__inst_mult_13_252 )))

	.dataa(!din_b[160]),
	.datab(!din_a[166]),
	.datac(!Xd_0__inst_mult_13_252 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_257 ),
	.sharein(Xd_0__inst_mult_13_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_177 ),
	.cout(Xd_0__inst_mult_13_178 ),
	.shareout(Xd_0__inst_mult_13_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_73 (
// Equation(s):
// Xd_0__inst_mult_15_192  = SUM(( !Xd_0__inst_mult_15_272  $ (((!din_b[184]) # (!din_a[190]))) ) + ( Xd_0__inst_mult_15_278  ) + ( Xd_0__inst_mult_15_277  ))
// Xd_0__inst_mult_15_193  = CARRY(( !Xd_0__inst_mult_15_272  $ (((!din_b[184]) # (!din_a[190]))) ) + ( Xd_0__inst_mult_15_278  ) + ( Xd_0__inst_mult_15_277  ))
// Xd_0__inst_mult_15_194  = SHARE((din_b[184] & (din_a[190] & Xd_0__inst_mult_15_272 )))

	.dataa(!din_b[184]),
	.datab(!din_a[190]),
	.datac(!Xd_0__inst_mult_15_272 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_277 ),
	.sharein(Xd_0__inst_mult_15_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_192 ),
	.cout(Xd_0__inst_mult_15_193 ),
	.shareout(Xd_0__inst_mult_15_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_68 (
// Equation(s):
// Xd_0__inst_mult_12_184  = SUM(( !Xd_0__inst_mult_12_264  $ (((!din_b[148]) # (!din_a[154]))) ) + ( Xd_0__inst_mult_12_270  ) + ( Xd_0__inst_mult_12_269  ))
// Xd_0__inst_mult_12_185  = CARRY(( !Xd_0__inst_mult_12_264  $ (((!din_b[148]) # (!din_a[154]))) ) + ( Xd_0__inst_mult_12_270  ) + ( Xd_0__inst_mult_12_269  ))
// Xd_0__inst_mult_12_186  = SHARE((din_b[148] & (din_a[154] & Xd_0__inst_mult_12_264 )))

	.dataa(!din_b[148]),
	.datab(!din_a[154]),
	.datac(!Xd_0__inst_mult_12_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_269 ),
	.sharein(Xd_0__inst_mult_12_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_184 ),
	.cout(Xd_0__inst_mult_12_185 ),
	.shareout(Xd_0__inst_mult_12_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_69 (
// Equation(s):
// Xd_0__inst_mult_12_188  = SUM(( (!din_a[151] & (((din_a[150] & din_b[154])))) # (din_a[151] & (!din_b[153] $ (((!din_a[150]) # (!din_b[154]))))) ) + ( Xd_0__inst_mult_12_274  ) + ( Xd_0__inst_mult_12_273  ))
// Xd_0__inst_mult_12_189  = CARRY(( (!din_a[151] & (((din_a[150] & din_b[154])))) # (din_a[151] & (!din_b[153] $ (((!din_a[150]) # (!din_b[154]))))) ) + ( Xd_0__inst_mult_12_274  ) + ( Xd_0__inst_mult_12_273  ))
// Xd_0__inst_mult_12_190  = SHARE((din_a[151] & (din_b[153] & (din_a[150] & din_b[154]))))

	.dataa(!din_a[151]),
	.datab(!din_b[153]),
	.datac(!din_a[150]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_273 ),
	.sharein(Xd_0__inst_mult_12_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_188 ),
	.cout(Xd_0__inst_mult_12_189 ),
	.shareout(Xd_0__inst_mult_12_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_73 (
// Equation(s):
// Xd_0__inst_mult_4_192  = SUM(( (din_a[53] & din_b[57]) ) + ( Xd_0__inst_mult_4_270  ) + ( Xd_0__inst_mult_4_269  ))
// Xd_0__inst_mult_4_193  = CARRY(( (din_a[53] & din_b[57]) ) + ( Xd_0__inst_mult_4_270  ) + ( Xd_0__inst_mult_4_269  ))
// Xd_0__inst_mult_4_194  = SHARE((din_a[53] & din_b[58]))

	.dataa(!din_a[53]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_269 ),
	.sharein(Xd_0__inst_mult_4_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_192 ),
	.cout(Xd_0__inst_mult_4_193 ),
	.shareout(Xd_0__inst_mult_4_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_70 (
// Equation(s):
// Xd_0__inst_mult_12_192  = SUM(( !Xd_0__inst_mult_12_0_q  $ (!Xd_0__inst_mult_12_1_q ) ) + ( Xd_0__inst_mult_12_37  ) + ( Xd_0__inst_mult_12_36  ))
// Xd_0__inst_mult_12_193  = CARRY(( !Xd_0__inst_mult_12_0_q  $ (!Xd_0__inst_mult_12_1_q ) ) + ( Xd_0__inst_mult_12_37  ) + ( Xd_0__inst_mult_12_36  ))
// Xd_0__inst_mult_12_194  = SHARE((Xd_0__inst_mult_12_0_q  & Xd_0__inst_mult_12_1_q ))

	.dataa(!Xd_0__inst_mult_12_0_q ),
	.datab(!Xd_0__inst_mult_12_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_36 ),
	.sharein(Xd_0__inst_mult_12_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_192 ),
	.cout(Xd_0__inst_mult_12_193 ),
	.shareout(Xd_0__inst_mult_12_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_70 (
// Equation(s):
// Xd_0__inst_mult_13_180  = SUM(( !Xd_0__inst_mult_13_0_q  $ (!Xd_0__inst_mult_13_1_q ) ) + ( Xd_0__inst_mult_1_37  ) + ( Xd_0__inst_mult_1_36  ))
// Xd_0__inst_mult_13_181  = CARRY(( !Xd_0__inst_mult_13_0_q  $ (!Xd_0__inst_mult_13_1_q ) ) + ( Xd_0__inst_mult_1_37  ) + ( Xd_0__inst_mult_1_36  ))
// Xd_0__inst_mult_13_182  = SHARE((Xd_0__inst_mult_13_0_q  & Xd_0__inst_mult_13_1_q ))

	.dataa(!Xd_0__inst_mult_13_0_q ),
	.datab(!Xd_0__inst_mult_13_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_36 ),
	.sharein(Xd_0__inst_mult_1_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_180 ),
	.cout(Xd_0__inst_mult_13_181 ),
	.shareout(Xd_0__inst_mult_13_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_74 (
// Equation(s):
// Xd_0__inst_mult_14_196  = SUM(( !Xd_0__inst_mult_14_0_q  $ (!Xd_0__inst_mult_14_1_q ) ) + ( Xd_0__inst_mult_6_37  ) + ( Xd_0__inst_mult_6_36  ))
// Xd_0__inst_mult_14_197  = CARRY(( !Xd_0__inst_mult_14_0_q  $ (!Xd_0__inst_mult_14_1_q ) ) + ( Xd_0__inst_mult_6_37  ) + ( Xd_0__inst_mult_6_36  ))
// Xd_0__inst_mult_14_198  = SHARE((Xd_0__inst_mult_14_0_q  & Xd_0__inst_mult_14_1_q ))

	.dataa(!Xd_0__inst_mult_14_0_q ),
	.datab(!Xd_0__inst_mult_14_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_36 ),
	.sharein(Xd_0__inst_mult_6_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_196 ),
	.cout(Xd_0__inst_mult_14_197 ),
	.shareout(Xd_0__inst_mult_14_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_74 (
// Equation(s):
// Xd_0__inst_mult_15_196  = SUM(( !Xd_0__inst_mult_15_0_q  $ (!Xd_0__inst_mult_15_1_q ) ) + ( Xd_0__inst_mult_5_37  ) + ( Xd_0__inst_mult_5_36  ))
// Xd_0__inst_mult_15_197  = CARRY(( !Xd_0__inst_mult_15_0_q  $ (!Xd_0__inst_mult_15_1_q ) ) + ( Xd_0__inst_mult_5_37  ) + ( Xd_0__inst_mult_5_36  ))
// Xd_0__inst_mult_15_198  = SHARE((Xd_0__inst_mult_15_0_q  & Xd_0__inst_mult_15_1_q ))

	.dataa(!Xd_0__inst_mult_15_0_q ),
	.datab(!Xd_0__inst_mult_15_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_36 ),
	.sharein(Xd_0__inst_mult_5_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_196 ),
	.cout(Xd_0__inst_mult_15_197 ),
	.shareout(Xd_0__inst_mult_15_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_66 (
// Equation(s):
// Xd_0__inst_mult_10_176  = SUM(( !Xd_0__inst_mult_10_0_q  $ (!Xd_0__inst_mult_10_1_q ) ) + ( Xd_0__inst_mult_2_37  ) + ( Xd_0__inst_mult_2_36  ))
// Xd_0__inst_mult_10_177  = CARRY(( !Xd_0__inst_mult_10_0_q  $ (!Xd_0__inst_mult_10_1_q ) ) + ( Xd_0__inst_mult_2_37  ) + ( Xd_0__inst_mult_2_36  ))
// Xd_0__inst_mult_10_178  = SHARE((Xd_0__inst_mult_10_0_q  & Xd_0__inst_mult_10_1_q ))

	.dataa(!Xd_0__inst_mult_10_0_q ),
	.datab(!Xd_0__inst_mult_10_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_36 ),
	.sharein(Xd_0__inst_mult_2_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_176 ),
	.cout(Xd_0__inst_mult_10_177 ),
	.shareout(Xd_0__inst_mult_10_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_70 (
// Equation(s):
// Xd_0__inst_mult_11_180  = SUM(( !Xd_0__inst_mult_11_0_q  $ (!Xd_0__inst_mult_11_1_q ) ) + ( Xd_0__inst_mult_14_37  ) + ( Xd_0__inst_mult_14_36  ))
// Xd_0__inst_mult_11_181  = CARRY(( !Xd_0__inst_mult_11_0_q  $ (!Xd_0__inst_mult_11_1_q ) ) + ( Xd_0__inst_mult_14_37  ) + ( Xd_0__inst_mult_14_36  ))
// Xd_0__inst_mult_11_182  = SHARE((Xd_0__inst_mult_11_0_q  & Xd_0__inst_mult_11_1_q ))

	.dataa(!Xd_0__inst_mult_11_0_q ),
	.datab(!Xd_0__inst_mult_11_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_36 ),
	.sharein(Xd_0__inst_mult_14_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_180 ),
	.cout(Xd_0__inst_mult_11_181 ),
	.shareout(Xd_0__inst_mult_11_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_70 (
// Equation(s):
// Xd_0__inst_mult_8_180  = SUM(( !Xd_0__inst_mult_8_0_q  $ (!Xd_0__inst_mult_8_1_q ) ) + ( Xd_0__inst_mult_12_41  ) + ( Xd_0__inst_mult_12_40  ))
// Xd_0__inst_mult_8_181  = CARRY(( !Xd_0__inst_mult_8_0_q  $ (!Xd_0__inst_mult_8_1_q ) ) + ( Xd_0__inst_mult_12_41  ) + ( Xd_0__inst_mult_12_40  ))
// Xd_0__inst_mult_8_182  = SHARE((Xd_0__inst_mult_8_0_q  & Xd_0__inst_mult_8_1_q ))

	.dataa(!Xd_0__inst_mult_8_0_q ),
	.datab(!Xd_0__inst_mult_8_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_40 ),
	.sharein(Xd_0__inst_mult_12_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_180 ),
	.cout(Xd_0__inst_mult_8_181 ),
	.shareout(Xd_0__inst_mult_8_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_66 (
// Equation(s):
// Xd_0__inst_mult_9_176  = SUM(( !Xd_0__inst_mult_9_0_q  $ (!Xd_0__inst_mult_9_1_q ) ) + ( Xd_0__inst_mult_15_37  ) + ( Xd_0__inst_mult_15_36  ))
// Xd_0__inst_mult_9_177  = CARRY(( !Xd_0__inst_mult_9_0_q  $ (!Xd_0__inst_mult_9_1_q ) ) + ( Xd_0__inst_mult_15_37  ) + ( Xd_0__inst_mult_15_36  ))
// Xd_0__inst_mult_9_178  = SHARE((Xd_0__inst_mult_9_0_q  & Xd_0__inst_mult_9_1_q ))

	.dataa(!Xd_0__inst_mult_9_0_q ),
	.datab(!Xd_0__inst_mult_9_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_36 ),
	.sharein(Xd_0__inst_mult_15_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_176 ),
	.cout(Xd_0__inst_mult_9_177 ),
	.shareout(Xd_0__inst_mult_9_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_66 (
// Equation(s):
// Xd_0__inst_mult_6_176  = SUM(( !Xd_0__inst_mult_6_0_q  $ (!Xd_0__inst_mult_6_1_q ) ) + ( Xd_0__inst_mult_5_41  ) + ( Xd_0__inst_mult_5_40  ))
// Xd_0__inst_mult_6_177  = CARRY(( !Xd_0__inst_mult_6_0_q  $ (!Xd_0__inst_mult_6_1_q ) ) + ( Xd_0__inst_mult_5_41  ) + ( Xd_0__inst_mult_5_40  ))
// Xd_0__inst_mult_6_178  = SHARE((Xd_0__inst_mult_6_0_q  & Xd_0__inst_mult_6_1_q ))

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_40 ),
	.sharein(Xd_0__inst_mult_5_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_176 ),
	.cout(Xd_0__inst_mult_6_177 ),
	.shareout(Xd_0__inst_mult_6_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_168 (
// Equation(s):
// Xd_0__inst_mult_7_169  = SUM(( !Xd_0__inst_mult_7_0_q  $ (!Xd_0__inst_mult_7_1_q ) ) + ( Xd_0__inst_mult_4_37  ) + ( Xd_0__inst_mult_4_36  ))
// Xd_0__inst_mult_7_170  = CARRY(( !Xd_0__inst_mult_7_0_q  $ (!Xd_0__inst_mult_7_1_q ) ) + ( Xd_0__inst_mult_4_37  ) + ( Xd_0__inst_mult_4_36  ))
// Xd_0__inst_mult_7_171  = SHARE((Xd_0__inst_mult_7_0_q  & Xd_0__inst_mult_7_1_q ))

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_36 ),
	.sharein(Xd_0__inst_mult_4_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_169 ),
	.cout(Xd_0__inst_mult_7_170 ),
	.shareout(Xd_0__inst_mult_7_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_74 (
// Equation(s):
// Xd_0__inst_mult_4_196  = SUM(( !Xd_0__inst_mult_4_0_q  $ (!Xd_0__inst_mult_4_1_q ) ) + ( Xd_0__inst_mult_10_37  ) + ( Xd_0__inst_mult_10_36  ))
// Xd_0__inst_mult_4_197  = CARRY(( !Xd_0__inst_mult_4_0_q  $ (!Xd_0__inst_mult_4_1_q ) ) + ( Xd_0__inst_mult_10_37  ) + ( Xd_0__inst_mult_10_36  ))
// Xd_0__inst_mult_4_198  = SHARE((Xd_0__inst_mult_4_0_q  & Xd_0__inst_mult_4_1_q ))

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_36 ),
	.sharein(Xd_0__inst_mult_10_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_196 ),
	.cout(Xd_0__inst_mult_4_197 ),
	.shareout(Xd_0__inst_mult_4_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_168 (
// Equation(s):
// Xd_0__inst_mult_5_169  = SUM(( !Xd_0__inst_mult_5_0_q  $ (!Xd_0__inst_mult_5_1_q ) ) + ( Xd_0__inst_mult_6_41  ) + ( Xd_0__inst_mult_6_40  ))
// Xd_0__inst_mult_5_170  = CARRY(( !Xd_0__inst_mult_5_0_q  $ (!Xd_0__inst_mult_5_1_q ) ) + ( Xd_0__inst_mult_6_41  ) + ( Xd_0__inst_mult_6_40  ))
// Xd_0__inst_mult_5_171  = SHARE((Xd_0__inst_mult_5_0_q  & Xd_0__inst_mult_5_1_q ))

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_40 ),
	.sharein(Xd_0__inst_mult_6_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_169 ),
	.cout(Xd_0__inst_mult_5_170 ),
	.shareout(Xd_0__inst_mult_5_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_172 (
// Equation(s):
// Xd_0__inst_mult_2_173  = SUM(( !Xd_0__inst_mult_2_0_q  $ (!Xd_0__inst_mult_2_1_q ) ) + ( Xd_0__inst_mult_2_41  ) + ( Xd_0__inst_mult_2_40  ))
// Xd_0__inst_mult_2_174  = CARRY(( !Xd_0__inst_mult_2_0_q  $ (!Xd_0__inst_mult_2_1_q ) ) + ( Xd_0__inst_mult_2_41  ) + ( Xd_0__inst_mult_2_40  ))
// Xd_0__inst_mult_2_175  = SHARE((Xd_0__inst_mult_2_0_q  & Xd_0__inst_mult_2_1_q ))

	.dataa(!Xd_0__inst_mult_2_0_q ),
	.datab(!Xd_0__inst_mult_2_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_40 ),
	.sharein(Xd_0__inst_mult_2_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_173 ),
	.cout(Xd_0__inst_mult_2_174 ),
	.shareout(Xd_0__inst_mult_2_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_168 (
// Equation(s):
// Xd_0__inst_mult_3_169  = SUM(( !Xd_0__inst_mult_3_0_q  $ (!Xd_0__inst_mult_3_1_q ) ) + ( Xd_0__inst_mult_13_37  ) + ( Xd_0__inst_mult_13_36  ))
// Xd_0__inst_mult_3_170  = CARRY(( !Xd_0__inst_mult_3_0_q  $ (!Xd_0__inst_mult_3_1_q ) ) + ( Xd_0__inst_mult_13_37  ) + ( Xd_0__inst_mult_13_36  ))
// Xd_0__inst_mult_3_171  = SHARE((Xd_0__inst_mult_3_0_q  & Xd_0__inst_mult_3_1_q ))

	.dataa(!Xd_0__inst_mult_3_0_q ),
	.datab(!Xd_0__inst_mult_3_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_36 ),
	.sharein(Xd_0__inst_mult_13_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_169 ),
	.cout(Xd_0__inst_mult_3_170 ),
	.shareout(Xd_0__inst_mult_3_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_172 (
// Equation(s):
// Xd_0__inst_mult_0_173  = SUM(( !Xd_0__inst_mult_0_0_q  $ (!Xd_0__inst_mult_0_1_q ) ) + ( Xd_0__inst_mult_14_41  ) + ( Xd_0__inst_mult_14_40  ))
// Xd_0__inst_mult_0_174  = CARRY(( !Xd_0__inst_mult_0_0_q  $ (!Xd_0__inst_mult_0_1_q ) ) + ( Xd_0__inst_mult_14_41  ) + ( Xd_0__inst_mult_14_40  ))
// Xd_0__inst_mult_0_175  = SHARE((Xd_0__inst_mult_0_0_q  & Xd_0__inst_mult_0_1_q ))

	.dataa(!Xd_0__inst_mult_0_0_q ),
	.datab(!Xd_0__inst_mult_0_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_40 ),
	.sharein(Xd_0__inst_mult_14_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_173 ),
	.cout(Xd_0__inst_mult_0_174 ),
	.shareout(Xd_0__inst_mult_0_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_172 (
// Equation(s):
// Xd_0__inst_mult_1_173  = SUM(( !Xd_0__inst_mult_1_0_q  $ (!Xd_0__inst_mult_1_1_q ) ) + ( Xd_0__inst_mult_3_37  ) + ( Xd_0__inst_mult_3_36  ))
// Xd_0__inst_mult_1_174  = CARRY(( !Xd_0__inst_mult_1_0_q  $ (!Xd_0__inst_mult_1_1_q ) ) + ( Xd_0__inst_mult_3_37  ) + ( Xd_0__inst_mult_3_36  ))
// Xd_0__inst_mult_1_175  = SHARE((Xd_0__inst_mult_1_0_q  & Xd_0__inst_mult_1_1_q ))

	.dataa(!Xd_0__inst_mult_1_0_q ),
	.datab(!Xd_0__inst_mult_1_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_36 ),
	.sharein(Xd_0__inst_mult_3_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_173 ),
	.cout(Xd_0__inst_mult_1_174 ),
	.shareout(Xd_0__inst_mult_1_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_71 (
// Equation(s):
// Xd_0__inst_mult_12_196  = SUM(( !Xd_0__inst_mult_12_2_q  $ (!Xd_0__inst_mult_12_3_q ) ) + ( Xd_0__inst_mult_12_194  ) + ( Xd_0__inst_mult_12_193  ))
// Xd_0__inst_mult_12_197  = CARRY(( !Xd_0__inst_mult_12_2_q  $ (!Xd_0__inst_mult_12_3_q ) ) + ( Xd_0__inst_mult_12_194  ) + ( Xd_0__inst_mult_12_193  ))
// Xd_0__inst_mult_12_198  = SHARE((Xd_0__inst_mult_12_2_q  & Xd_0__inst_mult_12_3_q ))

	.dataa(!Xd_0__inst_mult_12_2_q ),
	.datab(!Xd_0__inst_mult_12_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_193 ),
	.sharein(Xd_0__inst_mult_12_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_196 ),
	.cout(Xd_0__inst_mult_12_197 ),
	.shareout(Xd_0__inst_mult_12_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_71 (
// Equation(s):
// Xd_0__inst_mult_13_184  = SUM(( !Xd_0__inst_mult_13_2_q  $ (!Xd_0__inst_mult_13_3_q ) ) + ( Xd_0__inst_mult_13_182  ) + ( Xd_0__inst_mult_13_181  ))
// Xd_0__inst_mult_13_185  = CARRY(( !Xd_0__inst_mult_13_2_q  $ (!Xd_0__inst_mult_13_3_q ) ) + ( Xd_0__inst_mult_13_182  ) + ( Xd_0__inst_mult_13_181  ))
// Xd_0__inst_mult_13_186  = SHARE((Xd_0__inst_mult_13_2_q  & Xd_0__inst_mult_13_3_q ))

	.dataa(!Xd_0__inst_mult_13_2_q ),
	.datab(!Xd_0__inst_mult_13_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_181 ),
	.sharein(Xd_0__inst_mult_13_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_184 ),
	.cout(Xd_0__inst_mult_13_185 ),
	.shareout(Xd_0__inst_mult_13_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_75 (
// Equation(s):
// Xd_0__inst_mult_14_200  = SUM(( !Xd_0__inst_mult_14_2_q  $ (!Xd_0__inst_mult_14_3_q ) ) + ( Xd_0__inst_mult_14_198  ) + ( Xd_0__inst_mult_14_197  ))
// Xd_0__inst_mult_14_201  = CARRY(( !Xd_0__inst_mult_14_2_q  $ (!Xd_0__inst_mult_14_3_q ) ) + ( Xd_0__inst_mult_14_198  ) + ( Xd_0__inst_mult_14_197  ))
// Xd_0__inst_mult_14_202  = SHARE((Xd_0__inst_mult_14_2_q  & Xd_0__inst_mult_14_3_q ))

	.dataa(!Xd_0__inst_mult_14_2_q ),
	.datab(!Xd_0__inst_mult_14_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_197 ),
	.sharein(Xd_0__inst_mult_14_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_200 ),
	.cout(Xd_0__inst_mult_14_201 ),
	.shareout(Xd_0__inst_mult_14_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_75 (
// Equation(s):
// Xd_0__inst_mult_15_200  = SUM(( !Xd_0__inst_mult_15_2_q  $ (!Xd_0__inst_mult_15_3_q ) ) + ( Xd_0__inst_mult_15_198  ) + ( Xd_0__inst_mult_15_197  ))
// Xd_0__inst_mult_15_201  = CARRY(( !Xd_0__inst_mult_15_2_q  $ (!Xd_0__inst_mult_15_3_q ) ) + ( Xd_0__inst_mult_15_198  ) + ( Xd_0__inst_mult_15_197  ))
// Xd_0__inst_mult_15_202  = SHARE((Xd_0__inst_mult_15_2_q  & Xd_0__inst_mult_15_3_q ))

	.dataa(!Xd_0__inst_mult_15_2_q ),
	.datab(!Xd_0__inst_mult_15_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_197 ),
	.sharein(Xd_0__inst_mult_15_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_200 ),
	.cout(Xd_0__inst_mult_15_201 ),
	.shareout(Xd_0__inst_mult_15_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_67 (
// Equation(s):
// Xd_0__inst_mult_10_180  = SUM(( !Xd_0__inst_mult_10_2_q  $ (!Xd_0__inst_mult_10_3_q ) ) + ( Xd_0__inst_mult_10_178  ) + ( Xd_0__inst_mult_10_177  ))
// Xd_0__inst_mult_10_181  = CARRY(( !Xd_0__inst_mult_10_2_q  $ (!Xd_0__inst_mult_10_3_q ) ) + ( Xd_0__inst_mult_10_178  ) + ( Xd_0__inst_mult_10_177  ))
// Xd_0__inst_mult_10_182  = SHARE((Xd_0__inst_mult_10_2_q  & Xd_0__inst_mult_10_3_q ))

	.dataa(!Xd_0__inst_mult_10_2_q ),
	.datab(!Xd_0__inst_mult_10_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_177 ),
	.sharein(Xd_0__inst_mult_10_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_180 ),
	.cout(Xd_0__inst_mult_10_181 ),
	.shareout(Xd_0__inst_mult_10_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_71 (
// Equation(s):
// Xd_0__inst_mult_11_184  = SUM(( !Xd_0__inst_mult_11_2_q  $ (!Xd_0__inst_mult_11_3_q ) ) + ( Xd_0__inst_mult_11_182  ) + ( Xd_0__inst_mult_11_181  ))
// Xd_0__inst_mult_11_185  = CARRY(( !Xd_0__inst_mult_11_2_q  $ (!Xd_0__inst_mult_11_3_q ) ) + ( Xd_0__inst_mult_11_182  ) + ( Xd_0__inst_mult_11_181  ))
// Xd_0__inst_mult_11_186  = SHARE((Xd_0__inst_mult_11_2_q  & Xd_0__inst_mult_11_3_q ))

	.dataa(!Xd_0__inst_mult_11_2_q ),
	.datab(!Xd_0__inst_mult_11_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_181 ),
	.sharein(Xd_0__inst_mult_11_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_184 ),
	.cout(Xd_0__inst_mult_11_185 ),
	.shareout(Xd_0__inst_mult_11_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_71 (
// Equation(s):
// Xd_0__inst_mult_8_184  = SUM(( !Xd_0__inst_mult_8_2_q  $ (!Xd_0__inst_mult_8_3_q ) ) + ( Xd_0__inst_mult_8_182  ) + ( Xd_0__inst_mult_8_181  ))
// Xd_0__inst_mult_8_185  = CARRY(( !Xd_0__inst_mult_8_2_q  $ (!Xd_0__inst_mult_8_3_q ) ) + ( Xd_0__inst_mult_8_182  ) + ( Xd_0__inst_mult_8_181  ))
// Xd_0__inst_mult_8_186  = SHARE((Xd_0__inst_mult_8_2_q  & Xd_0__inst_mult_8_3_q ))

	.dataa(!Xd_0__inst_mult_8_2_q ),
	.datab(!Xd_0__inst_mult_8_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_181 ),
	.sharein(Xd_0__inst_mult_8_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_184 ),
	.cout(Xd_0__inst_mult_8_185 ),
	.shareout(Xd_0__inst_mult_8_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_67 (
// Equation(s):
// Xd_0__inst_mult_9_180  = SUM(( !Xd_0__inst_mult_9_2_q  $ (!Xd_0__inst_mult_9_3_q ) ) + ( Xd_0__inst_mult_9_178  ) + ( Xd_0__inst_mult_9_177  ))
// Xd_0__inst_mult_9_181  = CARRY(( !Xd_0__inst_mult_9_2_q  $ (!Xd_0__inst_mult_9_3_q ) ) + ( Xd_0__inst_mult_9_178  ) + ( Xd_0__inst_mult_9_177  ))
// Xd_0__inst_mult_9_182  = SHARE((Xd_0__inst_mult_9_2_q  & Xd_0__inst_mult_9_3_q ))

	.dataa(!Xd_0__inst_mult_9_2_q ),
	.datab(!Xd_0__inst_mult_9_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_177 ),
	.sharein(Xd_0__inst_mult_9_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_180 ),
	.cout(Xd_0__inst_mult_9_181 ),
	.shareout(Xd_0__inst_mult_9_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_67 (
// Equation(s):
// Xd_0__inst_mult_6_180  = SUM(( !Xd_0__inst_mult_6_2_q  $ (!Xd_0__inst_mult_6_3_q ) ) + ( Xd_0__inst_mult_6_178  ) + ( Xd_0__inst_mult_6_177  ))
// Xd_0__inst_mult_6_181  = CARRY(( !Xd_0__inst_mult_6_2_q  $ (!Xd_0__inst_mult_6_3_q ) ) + ( Xd_0__inst_mult_6_178  ) + ( Xd_0__inst_mult_6_177  ))
// Xd_0__inst_mult_6_182  = SHARE((Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_3_q ))

	.dataa(!Xd_0__inst_mult_6_2_q ),
	.datab(!Xd_0__inst_mult_6_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_177 ),
	.sharein(Xd_0__inst_mult_6_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_180 ),
	.cout(Xd_0__inst_mult_6_181 ),
	.shareout(Xd_0__inst_mult_6_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7 (
// Equation(s):
// Xd_0__inst_mult_7_173  = SUM(( !Xd_0__inst_mult_7_2_q  $ (!Xd_0__inst_mult_7_3_q ) ) + ( Xd_0__inst_mult_7_171  ) + ( Xd_0__inst_mult_7_170  ))
// Xd_0__inst_mult_7_174  = CARRY(( !Xd_0__inst_mult_7_2_q  $ (!Xd_0__inst_mult_7_3_q ) ) + ( Xd_0__inst_mult_7_171  ) + ( Xd_0__inst_mult_7_170  ))
// Xd_0__inst_mult_7_175  = SHARE((Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_3_q ))

	.dataa(!Xd_0__inst_mult_7_2_q ),
	.datab(!Xd_0__inst_mult_7_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_170 ),
	.sharein(Xd_0__inst_mult_7_171 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_173 ),
	.cout(Xd_0__inst_mult_7_174 ),
	.shareout(Xd_0__inst_mult_7_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_75 (
// Equation(s):
// Xd_0__inst_mult_4_200  = SUM(( !Xd_0__inst_mult_4_2_q  $ (!Xd_0__inst_mult_4_3_q ) ) + ( Xd_0__inst_mult_4_198  ) + ( Xd_0__inst_mult_4_197  ))
// Xd_0__inst_mult_4_201  = CARRY(( !Xd_0__inst_mult_4_2_q  $ (!Xd_0__inst_mult_4_3_q ) ) + ( Xd_0__inst_mult_4_198  ) + ( Xd_0__inst_mult_4_197  ))
// Xd_0__inst_mult_4_202  = SHARE((Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_3_q ))

	.dataa(!Xd_0__inst_mult_4_2_q ),
	.datab(!Xd_0__inst_mult_4_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_197 ),
	.sharein(Xd_0__inst_mult_4_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_200 ),
	.cout(Xd_0__inst_mult_4_201 ),
	.shareout(Xd_0__inst_mult_4_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5 (
// Equation(s):
// Xd_0__inst_mult_5_173  = SUM(( !Xd_0__inst_mult_5_2_q  $ (!Xd_0__inst_mult_5_3_q ) ) + ( Xd_0__inst_mult_5_171  ) + ( Xd_0__inst_mult_5_170  ))
// Xd_0__inst_mult_5_174  = CARRY(( !Xd_0__inst_mult_5_2_q  $ (!Xd_0__inst_mult_5_3_q ) ) + ( Xd_0__inst_mult_5_171  ) + ( Xd_0__inst_mult_5_170  ))
// Xd_0__inst_mult_5_175  = SHARE((Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_3_q ))

	.dataa(!Xd_0__inst_mult_5_2_q ),
	.datab(!Xd_0__inst_mult_5_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_170 ),
	.sharein(Xd_0__inst_mult_5_171 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_173 ),
	.cout(Xd_0__inst_mult_5_174 ),
	.shareout(Xd_0__inst_mult_5_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2 (
// Equation(s):
// Xd_0__inst_mult_2_177  = SUM(( !Xd_0__inst_mult_2_2_q  $ (!Xd_0__inst_mult_2_3_q ) ) + ( Xd_0__inst_mult_2_175  ) + ( Xd_0__inst_mult_2_174  ))
// Xd_0__inst_mult_2_178  = CARRY(( !Xd_0__inst_mult_2_2_q  $ (!Xd_0__inst_mult_2_3_q ) ) + ( Xd_0__inst_mult_2_175  ) + ( Xd_0__inst_mult_2_174  ))
// Xd_0__inst_mult_2_179  = SHARE((Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_3_q ))

	.dataa(!Xd_0__inst_mult_2_2_q ),
	.datab(!Xd_0__inst_mult_2_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_174 ),
	.sharein(Xd_0__inst_mult_2_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_177 ),
	.cout(Xd_0__inst_mult_2_178 ),
	.shareout(Xd_0__inst_mult_2_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3 (
// Equation(s):
// Xd_0__inst_mult_3_173  = SUM(( !Xd_0__inst_mult_3_2_q  $ (!Xd_0__inst_mult_3_3_q ) ) + ( Xd_0__inst_mult_3_171  ) + ( Xd_0__inst_mult_3_170  ))
// Xd_0__inst_mult_3_174  = CARRY(( !Xd_0__inst_mult_3_2_q  $ (!Xd_0__inst_mult_3_3_q ) ) + ( Xd_0__inst_mult_3_171  ) + ( Xd_0__inst_mult_3_170  ))
// Xd_0__inst_mult_3_175  = SHARE((Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_3_q ))

	.dataa(!Xd_0__inst_mult_3_2_q ),
	.datab(!Xd_0__inst_mult_3_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_170 ),
	.sharein(Xd_0__inst_mult_3_171 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_173 ),
	.cout(Xd_0__inst_mult_3_174 ),
	.shareout(Xd_0__inst_mult_3_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0 (
// Equation(s):
// Xd_0__inst_mult_0_177  = SUM(( !Xd_0__inst_mult_0_2_q  $ (!Xd_0__inst_mult_0_3_q ) ) + ( Xd_0__inst_mult_0_175  ) + ( Xd_0__inst_mult_0_174  ))
// Xd_0__inst_mult_0_178  = CARRY(( !Xd_0__inst_mult_0_2_q  $ (!Xd_0__inst_mult_0_3_q ) ) + ( Xd_0__inst_mult_0_175  ) + ( Xd_0__inst_mult_0_174  ))
// Xd_0__inst_mult_0_179  = SHARE((Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_3_q ))

	.dataa(!Xd_0__inst_mult_0_2_q ),
	.datab(!Xd_0__inst_mult_0_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_174 ),
	.sharein(Xd_0__inst_mult_0_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_177 ),
	.cout(Xd_0__inst_mult_0_178 ),
	.shareout(Xd_0__inst_mult_0_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1 (
// Equation(s):
// Xd_0__inst_mult_1_177  = SUM(( !Xd_0__inst_mult_1_2_q  $ (!Xd_0__inst_mult_1_3_q ) ) + ( Xd_0__inst_mult_1_175  ) + ( Xd_0__inst_mult_1_174  ))
// Xd_0__inst_mult_1_178  = CARRY(( !Xd_0__inst_mult_1_2_q  $ (!Xd_0__inst_mult_1_3_q ) ) + ( Xd_0__inst_mult_1_175  ) + ( Xd_0__inst_mult_1_174  ))
// Xd_0__inst_mult_1_179  = SHARE((Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_3_q ))

	.dataa(!Xd_0__inst_mult_1_2_q ),
	.datab(!Xd_0__inst_mult_1_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_174 ),
	.sharein(Xd_0__inst_mult_1_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_177 ),
	.cout(Xd_0__inst_mult_1_178 ),
	.shareout(Xd_0__inst_mult_1_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_72 (
// Equation(s):
// Xd_0__inst_mult_12_200  = SUM(( !Xd_0__inst_mult_12_4_q  $ (!Xd_0__inst_mult_12_5_q ) ) + ( Xd_0__inst_mult_12_198  ) + ( Xd_0__inst_mult_12_197  ))
// Xd_0__inst_mult_12_201  = CARRY(( !Xd_0__inst_mult_12_4_q  $ (!Xd_0__inst_mult_12_5_q ) ) + ( Xd_0__inst_mult_12_198  ) + ( Xd_0__inst_mult_12_197  ))
// Xd_0__inst_mult_12_202  = SHARE((Xd_0__inst_mult_12_4_q  & Xd_0__inst_mult_12_5_q ))

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_197 ),
	.sharein(Xd_0__inst_mult_12_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_200 ),
	.cout(Xd_0__inst_mult_12_201 ),
	.shareout(Xd_0__inst_mult_12_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_72 (
// Equation(s):
// Xd_0__inst_mult_13_188  = SUM(( !Xd_0__inst_mult_13_4_q  $ (!Xd_0__inst_mult_13_5_q ) ) + ( Xd_0__inst_mult_13_186  ) + ( Xd_0__inst_mult_13_185  ))
// Xd_0__inst_mult_13_189  = CARRY(( !Xd_0__inst_mult_13_4_q  $ (!Xd_0__inst_mult_13_5_q ) ) + ( Xd_0__inst_mult_13_186  ) + ( Xd_0__inst_mult_13_185  ))
// Xd_0__inst_mult_13_190  = SHARE((Xd_0__inst_mult_13_4_q  & Xd_0__inst_mult_13_5_q ))

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_185 ),
	.sharein(Xd_0__inst_mult_13_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_188 ),
	.cout(Xd_0__inst_mult_13_189 ),
	.shareout(Xd_0__inst_mult_13_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_76 (
// Equation(s):
// Xd_0__inst_mult_14_204  = SUM(( !Xd_0__inst_mult_14_4_q  $ (!Xd_0__inst_mult_14_5_q ) ) + ( Xd_0__inst_mult_14_202  ) + ( Xd_0__inst_mult_14_201  ))
// Xd_0__inst_mult_14_205  = CARRY(( !Xd_0__inst_mult_14_4_q  $ (!Xd_0__inst_mult_14_5_q ) ) + ( Xd_0__inst_mult_14_202  ) + ( Xd_0__inst_mult_14_201  ))
// Xd_0__inst_mult_14_206  = SHARE((Xd_0__inst_mult_14_4_q  & Xd_0__inst_mult_14_5_q ))

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_201 ),
	.sharein(Xd_0__inst_mult_14_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_204 ),
	.cout(Xd_0__inst_mult_14_205 ),
	.shareout(Xd_0__inst_mult_14_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_76 (
// Equation(s):
// Xd_0__inst_mult_15_204  = SUM(( !Xd_0__inst_mult_15_4_q  $ (!Xd_0__inst_mult_15_5_q ) ) + ( Xd_0__inst_mult_15_202  ) + ( Xd_0__inst_mult_15_201  ))
// Xd_0__inst_mult_15_205  = CARRY(( !Xd_0__inst_mult_15_4_q  $ (!Xd_0__inst_mult_15_5_q ) ) + ( Xd_0__inst_mult_15_202  ) + ( Xd_0__inst_mult_15_201  ))
// Xd_0__inst_mult_15_206  = SHARE((Xd_0__inst_mult_15_4_q  & Xd_0__inst_mult_15_5_q ))

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_201 ),
	.sharein(Xd_0__inst_mult_15_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_204 ),
	.cout(Xd_0__inst_mult_15_205 ),
	.shareout(Xd_0__inst_mult_15_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_68 (
// Equation(s):
// Xd_0__inst_mult_10_184  = SUM(( !Xd_0__inst_mult_10_4_q  $ (!Xd_0__inst_mult_10_5_q ) ) + ( Xd_0__inst_mult_10_182  ) + ( Xd_0__inst_mult_10_181  ))
// Xd_0__inst_mult_10_185  = CARRY(( !Xd_0__inst_mult_10_4_q  $ (!Xd_0__inst_mult_10_5_q ) ) + ( Xd_0__inst_mult_10_182  ) + ( Xd_0__inst_mult_10_181  ))
// Xd_0__inst_mult_10_186  = SHARE((Xd_0__inst_mult_10_4_q  & Xd_0__inst_mult_10_5_q ))

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_181 ),
	.sharein(Xd_0__inst_mult_10_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_184 ),
	.cout(Xd_0__inst_mult_10_185 ),
	.shareout(Xd_0__inst_mult_10_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_72 (
// Equation(s):
// Xd_0__inst_mult_11_188  = SUM(( !Xd_0__inst_mult_11_4_q  $ (!Xd_0__inst_mult_11_5_q ) ) + ( Xd_0__inst_mult_11_186  ) + ( Xd_0__inst_mult_11_185  ))
// Xd_0__inst_mult_11_189  = CARRY(( !Xd_0__inst_mult_11_4_q  $ (!Xd_0__inst_mult_11_5_q ) ) + ( Xd_0__inst_mult_11_186  ) + ( Xd_0__inst_mult_11_185  ))
// Xd_0__inst_mult_11_190  = SHARE((Xd_0__inst_mult_11_4_q  & Xd_0__inst_mult_11_5_q ))

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_185 ),
	.sharein(Xd_0__inst_mult_11_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_188 ),
	.cout(Xd_0__inst_mult_11_189 ),
	.shareout(Xd_0__inst_mult_11_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_72 (
// Equation(s):
// Xd_0__inst_mult_8_188  = SUM(( !Xd_0__inst_mult_8_4_q  $ (!Xd_0__inst_mult_8_5_q ) ) + ( Xd_0__inst_mult_8_186  ) + ( Xd_0__inst_mult_8_185  ))
// Xd_0__inst_mult_8_189  = CARRY(( !Xd_0__inst_mult_8_4_q  $ (!Xd_0__inst_mult_8_5_q ) ) + ( Xd_0__inst_mult_8_186  ) + ( Xd_0__inst_mult_8_185  ))
// Xd_0__inst_mult_8_190  = SHARE((Xd_0__inst_mult_8_4_q  & Xd_0__inst_mult_8_5_q ))

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_185 ),
	.sharein(Xd_0__inst_mult_8_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_188 ),
	.cout(Xd_0__inst_mult_8_189 ),
	.shareout(Xd_0__inst_mult_8_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_68 (
// Equation(s):
// Xd_0__inst_mult_9_184  = SUM(( !Xd_0__inst_mult_9_4_q  $ (!Xd_0__inst_mult_9_5_q ) ) + ( Xd_0__inst_mult_9_182  ) + ( Xd_0__inst_mult_9_181  ))
// Xd_0__inst_mult_9_185  = CARRY(( !Xd_0__inst_mult_9_4_q  $ (!Xd_0__inst_mult_9_5_q ) ) + ( Xd_0__inst_mult_9_182  ) + ( Xd_0__inst_mult_9_181  ))
// Xd_0__inst_mult_9_186  = SHARE((Xd_0__inst_mult_9_4_q  & Xd_0__inst_mult_9_5_q ))

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_181 ),
	.sharein(Xd_0__inst_mult_9_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_184 ),
	.cout(Xd_0__inst_mult_9_185 ),
	.shareout(Xd_0__inst_mult_9_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_68 (
// Equation(s):
// Xd_0__inst_mult_6_184  = SUM(( !Xd_0__inst_mult_6_4_q  $ (!Xd_0__inst_mult_6_5_q ) ) + ( Xd_0__inst_mult_6_182  ) + ( Xd_0__inst_mult_6_181  ))
// Xd_0__inst_mult_6_185  = CARRY(( !Xd_0__inst_mult_6_4_q  $ (!Xd_0__inst_mult_6_5_q ) ) + ( Xd_0__inst_mult_6_182  ) + ( Xd_0__inst_mult_6_181  ))
// Xd_0__inst_mult_6_186  = SHARE((Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_5_q ))

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_181 ),
	.sharein(Xd_0__inst_mult_6_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_184 ),
	.cout(Xd_0__inst_mult_6_185 ),
	.shareout(Xd_0__inst_mult_6_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_66 (
// Equation(s):
// Xd_0__inst_mult_7_176  = SUM(( !Xd_0__inst_mult_7_4_q  $ (!Xd_0__inst_mult_7_5_q ) ) + ( Xd_0__inst_mult_7_175  ) + ( Xd_0__inst_mult_7_174  ))
// Xd_0__inst_mult_7_177  = CARRY(( !Xd_0__inst_mult_7_4_q  $ (!Xd_0__inst_mult_7_5_q ) ) + ( Xd_0__inst_mult_7_175  ) + ( Xd_0__inst_mult_7_174  ))
// Xd_0__inst_mult_7_178  = SHARE((Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_5_q ))

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_174 ),
	.sharein(Xd_0__inst_mult_7_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_176 ),
	.cout(Xd_0__inst_mult_7_177 ),
	.shareout(Xd_0__inst_mult_7_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_76 (
// Equation(s):
// Xd_0__inst_mult_4_204  = SUM(( !Xd_0__inst_mult_4_4_q  $ (!Xd_0__inst_mult_4_5_q ) ) + ( Xd_0__inst_mult_4_202  ) + ( Xd_0__inst_mult_4_201  ))
// Xd_0__inst_mult_4_205  = CARRY(( !Xd_0__inst_mult_4_4_q  $ (!Xd_0__inst_mult_4_5_q ) ) + ( Xd_0__inst_mult_4_202  ) + ( Xd_0__inst_mult_4_201  ))
// Xd_0__inst_mult_4_206  = SHARE((Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_5_q ))

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_201 ),
	.sharein(Xd_0__inst_mult_4_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_204 ),
	.cout(Xd_0__inst_mult_4_205 ),
	.shareout(Xd_0__inst_mult_4_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_66 (
// Equation(s):
// Xd_0__inst_mult_5_176  = SUM(( !Xd_0__inst_mult_5_4_q  $ (!Xd_0__inst_mult_5_5_q ) ) + ( Xd_0__inst_mult_5_175  ) + ( Xd_0__inst_mult_5_174  ))
// Xd_0__inst_mult_5_177  = CARRY(( !Xd_0__inst_mult_5_4_q  $ (!Xd_0__inst_mult_5_5_q ) ) + ( Xd_0__inst_mult_5_175  ) + ( Xd_0__inst_mult_5_174  ))
// Xd_0__inst_mult_5_178  = SHARE((Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_5_q ))

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_174 ),
	.sharein(Xd_0__inst_mult_5_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_176 ),
	.cout(Xd_0__inst_mult_5_177 ),
	.shareout(Xd_0__inst_mult_5_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_70 (
// Equation(s):
// Xd_0__inst_mult_2_180  = SUM(( !Xd_0__inst_mult_2_4_q  $ (!Xd_0__inst_mult_2_5_q ) ) + ( Xd_0__inst_mult_2_179  ) + ( Xd_0__inst_mult_2_178  ))
// Xd_0__inst_mult_2_181  = CARRY(( !Xd_0__inst_mult_2_4_q  $ (!Xd_0__inst_mult_2_5_q ) ) + ( Xd_0__inst_mult_2_179  ) + ( Xd_0__inst_mult_2_178  ))
// Xd_0__inst_mult_2_182  = SHARE((Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_5_q ))

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_178 ),
	.sharein(Xd_0__inst_mult_2_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_180 ),
	.cout(Xd_0__inst_mult_2_181 ),
	.shareout(Xd_0__inst_mult_2_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_66 (
// Equation(s):
// Xd_0__inst_mult_3_176  = SUM(( !Xd_0__inst_mult_3_4_q  $ (!Xd_0__inst_mult_3_5_q ) ) + ( Xd_0__inst_mult_3_175  ) + ( Xd_0__inst_mult_3_174  ))
// Xd_0__inst_mult_3_177  = CARRY(( !Xd_0__inst_mult_3_4_q  $ (!Xd_0__inst_mult_3_5_q ) ) + ( Xd_0__inst_mult_3_175  ) + ( Xd_0__inst_mult_3_174  ))
// Xd_0__inst_mult_3_178  = SHARE((Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_5_q ))

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_174 ),
	.sharein(Xd_0__inst_mult_3_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_176 ),
	.cout(Xd_0__inst_mult_3_177 ),
	.shareout(Xd_0__inst_mult_3_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_70 (
// Equation(s):
// Xd_0__inst_mult_0_180  = SUM(( !Xd_0__inst_mult_0_4_q  $ (!Xd_0__inst_mult_0_5_q ) ) + ( Xd_0__inst_mult_0_179  ) + ( Xd_0__inst_mult_0_178  ))
// Xd_0__inst_mult_0_181  = CARRY(( !Xd_0__inst_mult_0_4_q  $ (!Xd_0__inst_mult_0_5_q ) ) + ( Xd_0__inst_mult_0_179  ) + ( Xd_0__inst_mult_0_178  ))
// Xd_0__inst_mult_0_182  = SHARE((Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_5_q ))

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_178 ),
	.sharein(Xd_0__inst_mult_0_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_180 ),
	.cout(Xd_0__inst_mult_0_181 ),
	.shareout(Xd_0__inst_mult_0_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_70 (
// Equation(s):
// Xd_0__inst_mult_1_180  = SUM(( !Xd_0__inst_mult_1_4_q  $ (!Xd_0__inst_mult_1_5_q ) ) + ( Xd_0__inst_mult_1_179  ) + ( Xd_0__inst_mult_1_178  ))
// Xd_0__inst_mult_1_181  = CARRY(( !Xd_0__inst_mult_1_4_q  $ (!Xd_0__inst_mult_1_5_q ) ) + ( Xd_0__inst_mult_1_179  ) + ( Xd_0__inst_mult_1_178  ))
// Xd_0__inst_mult_1_182  = SHARE((Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_5_q ))

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_178 ),
	.sharein(Xd_0__inst_mult_1_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_180 ),
	.cout(Xd_0__inst_mult_1_181 ),
	.shareout(Xd_0__inst_mult_1_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_73 (
// Equation(s):
// Xd_0__inst_mult_12_204  = SUM(( !Xd_0__inst_mult_12_6_q  $ (!Xd_0__inst_mult_12_7_q ) ) + ( Xd_0__inst_mult_12_202  ) + ( Xd_0__inst_mult_12_201  ))
// Xd_0__inst_mult_12_205  = CARRY(( !Xd_0__inst_mult_12_6_q  $ (!Xd_0__inst_mult_12_7_q ) ) + ( Xd_0__inst_mult_12_202  ) + ( Xd_0__inst_mult_12_201  ))
// Xd_0__inst_mult_12_206  = SHARE((Xd_0__inst_mult_12_6_q  & Xd_0__inst_mult_12_7_q ))

	.dataa(!Xd_0__inst_mult_12_6_q ),
	.datab(!Xd_0__inst_mult_12_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_201 ),
	.sharein(Xd_0__inst_mult_12_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_204 ),
	.cout(Xd_0__inst_mult_12_205 ),
	.shareout(Xd_0__inst_mult_12_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_73 (
// Equation(s):
// Xd_0__inst_mult_13_192  = SUM(( !Xd_0__inst_mult_13_6_q  $ (!Xd_0__inst_mult_13_7_q ) ) + ( Xd_0__inst_mult_13_190  ) + ( Xd_0__inst_mult_13_189  ))
// Xd_0__inst_mult_13_193  = CARRY(( !Xd_0__inst_mult_13_6_q  $ (!Xd_0__inst_mult_13_7_q ) ) + ( Xd_0__inst_mult_13_190  ) + ( Xd_0__inst_mult_13_189  ))
// Xd_0__inst_mult_13_194  = SHARE((Xd_0__inst_mult_13_6_q  & Xd_0__inst_mult_13_7_q ))

	.dataa(!Xd_0__inst_mult_13_6_q ),
	.datab(!Xd_0__inst_mult_13_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_189 ),
	.sharein(Xd_0__inst_mult_13_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_192 ),
	.cout(Xd_0__inst_mult_13_193 ),
	.shareout(Xd_0__inst_mult_13_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_77 (
// Equation(s):
// Xd_0__inst_mult_14_208  = SUM(( !Xd_0__inst_mult_14_6_q  $ (!Xd_0__inst_mult_14_7_q ) ) + ( Xd_0__inst_mult_14_206  ) + ( Xd_0__inst_mult_14_205  ))
// Xd_0__inst_mult_14_209  = CARRY(( !Xd_0__inst_mult_14_6_q  $ (!Xd_0__inst_mult_14_7_q ) ) + ( Xd_0__inst_mult_14_206  ) + ( Xd_0__inst_mult_14_205  ))
// Xd_0__inst_mult_14_210  = SHARE((Xd_0__inst_mult_14_6_q  & Xd_0__inst_mult_14_7_q ))

	.dataa(!Xd_0__inst_mult_14_6_q ),
	.datab(!Xd_0__inst_mult_14_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_205 ),
	.sharein(Xd_0__inst_mult_14_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_208 ),
	.cout(Xd_0__inst_mult_14_209 ),
	.shareout(Xd_0__inst_mult_14_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_77 (
// Equation(s):
// Xd_0__inst_mult_15_208  = SUM(( !Xd_0__inst_mult_15_6_q  $ (!Xd_0__inst_mult_15_7_q ) ) + ( Xd_0__inst_mult_15_206  ) + ( Xd_0__inst_mult_15_205  ))
// Xd_0__inst_mult_15_209  = CARRY(( !Xd_0__inst_mult_15_6_q  $ (!Xd_0__inst_mult_15_7_q ) ) + ( Xd_0__inst_mult_15_206  ) + ( Xd_0__inst_mult_15_205  ))
// Xd_0__inst_mult_15_210  = SHARE((Xd_0__inst_mult_15_6_q  & Xd_0__inst_mult_15_7_q ))

	.dataa(!Xd_0__inst_mult_15_6_q ),
	.datab(!Xd_0__inst_mult_15_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_205 ),
	.sharein(Xd_0__inst_mult_15_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_208 ),
	.cout(Xd_0__inst_mult_15_209 ),
	.shareout(Xd_0__inst_mult_15_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_69 (
// Equation(s):
// Xd_0__inst_mult_10_188  = SUM(( !Xd_0__inst_mult_10_6_q  $ (!Xd_0__inst_mult_10_7_q ) ) + ( Xd_0__inst_mult_10_186  ) + ( Xd_0__inst_mult_10_185  ))
// Xd_0__inst_mult_10_189  = CARRY(( !Xd_0__inst_mult_10_6_q  $ (!Xd_0__inst_mult_10_7_q ) ) + ( Xd_0__inst_mult_10_186  ) + ( Xd_0__inst_mult_10_185  ))
// Xd_0__inst_mult_10_190  = SHARE((Xd_0__inst_mult_10_6_q  & Xd_0__inst_mult_10_7_q ))

	.dataa(!Xd_0__inst_mult_10_6_q ),
	.datab(!Xd_0__inst_mult_10_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_185 ),
	.sharein(Xd_0__inst_mult_10_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_188 ),
	.cout(Xd_0__inst_mult_10_189 ),
	.shareout(Xd_0__inst_mult_10_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_73 (
// Equation(s):
// Xd_0__inst_mult_11_192  = SUM(( !Xd_0__inst_mult_11_6_q  $ (!Xd_0__inst_mult_11_7_q ) ) + ( Xd_0__inst_mult_11_190  ) + ( Xd_0__inst_mult_11_189  ))
// Xd_0__inst_mult_11_193  = CARRY(( !Xd_0__inst_mult_11_6_q  $ (!Xd_0__inst_mult_11_7_q ) ) + ( Xd_0__inst_mult_11_190  ) + ( Xd_0__inst_mult_11_189  ))
// Xd_0__inst_mult_11_194  = SHARE((Xd_0__inst_mult_11_6_q  & Xd_0__inst_mult_11_7_q ))

	.dataa(!Xd_0__inst_mult_11_6_q ),
	.datab(!Xd_0__inst_mult_11_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_189 ),
	.sharein(Xd_0__inst_mult_11_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_192 ),
	.cout(Xd_0__inst_mult_11_193 ),
	.shareout(Xd_0__inst_mult_11_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_73 (
// Equation(s):
// Xd_0__inst_mult_8_192  = SUM(( !Xd_0__inst_mult_8_6_q  $ (!Xd_0__inst_mult_8_7_q ) ) + ( Xd_0__inst_mult_8_190  ) + ( Xd_0__inst_mult_8_189  ))
// Xd_0__inst_mult_8_193  = CARRY(( !Xd_0__inst_mult_8_6_q  $ (!Xd_0__inst_mult_8_7_q ) ) + ( Xd_0__inst_mult_8_190  ) + ( Xd_0__inst_mult_8_189  ))
// Xd_0__inst_mult_8_194  = SHARE((Xd_0__inst_mult_8_6_q  & Xd_0__inst_mult_8_7_q ))

	.dataa(!Xd_0__inst_mult_8_6_q ),
	.datab(!Xd_0__inst_mult_8_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_189 ),
	.sharein(Xd_0__inst_mult_8_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_192 ),
	.cout(Xd_0__inst_mult_8_193 ),
	.shareout(Xd_0__inst_mult_8_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_69 (
// Equation(s):
// Xd_0__inst_mult_9_188  = SUM(( !Xd_0__inst_mult_9_6_q  $ (!Xd_0__inst_mult_9_7_q ) ) + ( Xd_0__inst_mult_9_186  ) + ( Xd_0__inst_mult_9_185  ))
// Xd_0__inst_mult_9_189  = CARRY(( !Xd_0__inst_mult_9_6_q  $ (!Xd_0__inst_mult_9_7_q ) ) + ( Xd_0__inst_mult_9_186  ) + ( Xd_0__inst_mult_9_185  ))
// Xd_0__inst_mult_9_190  = SHARE((Xd_0__inst_mult_9_6_q  & Xd_0__inst_mult_9_7_q ))

	.dataa(!Xd_0__inst_mult_9_6_q ),
	.datab(!Xd_0__inst_mult_9_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_185 ),
	.sharein(Xd_0__inst_mult_9_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_188 ),
	.cout(Xd_0__inst_mult_9_189 ),
	.shareout(Xd_0__inst_mult_9_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_69 (
// Equation(s):
// Xd_0__inst_mult_6_188  = SUM(( !Xd_0__inst_mult_6_6_q  $ (!Xd_0__inst_mult_6_7_q ) ) + ( Xd_0__inst_mult_6_186  ) + ( Xd_0__inst_mult_6_185  ))
// Xd_0__inst_mult_6_189  = CARRY(( !Xd_0__inst_mult_6_6_q  $ (!Xd_0__inst_mult_6_7_q ) ) + ( Xd_0__inst_mult_6_186  ) + ( Xd_0__inst_mult_6_185  ))
// Xd_0__inst_mult_6_190  = SHARE((Xd_0__inst_mult_6_6_q  & Xd_0__inst_mult_6_7_q ))

	.dataa(!Xd_0__inst_mult_6_6_q ),
	.datab(!Xd_0__inst_mult_6_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_185 ),
	.sharein(Xd_0__inst_mult_6_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_188 ),
	.cout(Xd_0__inst_mult_6_189 ),
	.shareout(Xd_0__inst_mult_6_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_67 (
// Equation(s):
// Xd_0__inst_mult_7_180  = SUM(( !Xd_0__inst_mult_7_6_q  $ (!Xd_0__inst_mult_7_7_q ) ) + ( Xd_0__inst_mult_7_178  ) + ( Xd_0__inst_mult_7_177  ))
// Xd_0__inst_mult_7_181  = CARRY(( !Xd_0__inst_mult_7_6_q  $ (!Xd_0__inst_mult_7_7_q ) ) + ( Xd_0__inst_mult_7_178  ) + ( Xd_0__inst_mult_7_177  ))
// Xd_0__inst_mult_7_182  = SHARE((Xd_0__inst_mult_7_6_q  & Xd_0__inst_mult_7_7_q ))

	.dataa(!Xd_0__inst_mult_7_6_q ),
	.datab(!Xd_0__inst_mult_7_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_177 ),
	.sharein(Xd_0__inst_mult_7_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_180 ),
	.cout(Xd_0__inst_mult_7_181 ),
	.shareout(Xd_0__inst_mult_7_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_77 (
// Equation(s):
// Xd_0__inst_mult_4_208  = SUM(( !Xd_0__inst_mult_4_6_q  $ (!Xd_0__inst_mult_4_7_q ) ) + ( Xd_0__inst_mult_4_206  ) + ( Xd_0__inst_mult_4_205  ))
// Xd_0__inst_mult_4_209  = CARRY(( !Xd_0__inst_mult_4_6_q  $ (!Xd_0__inst_mult_4_7_q ) ) + ( Xd_0__inst_mult_4_206  ) + ( Xd_0__inst_mult_4_205  ))
// Xd_0__inst_mult_4_210  = SHARE((Xd_0__inst_mult_4_6_q  & Xd_0__inst_mult_4_7_q ))

	.dataa(!Xd_0__inst_mult_4_6_q ),
	.datab(!Xd_0__inst_mult_4_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_205 ),
	.sharein(Xd_0__inst_mult_4_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_208 ),
	.cout(Xd_0__inst_mult_4_209 ),
	.shareout(Xd_0__inst_mult_4_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_67 (
// Equation(s):
// Xd_0__inst_mult_5_180  = SUM(( !Xd_0__inst_mult_5_6_q  $ (!Xd_0__inst_mult_5_7_q ) ) + ( Xd_0__inst_mult_5_178  ) + ( Xd_0__inst_mult_5_177  ))
// Xd_0__inst_mult_5_181  = CARRY(( !Xd_0__inst_mult_5_6_q  $ (!Xd_0__inst_mult_5_7_q ) ) + ( Xd_0__inst_mult_5_178  ) + ( Xd_0__inst_mult_5_177  ))
// Xd_0__inst_mult_5_182  = SHARE((Xd_0__inst_mult_5_6_q  & Xd_0__inst_mult_5_7_q ))

	.dataa(!Xd_0__inst_mult_5_6_q ),
	.datab(!Xd_0__inst_mult_5_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_177 ),
	.sharein(Xd_0__inst_mult_5_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_180 ),
	.cout(Xd_0__inst_mult_5_181 ),
	.shareout(Xd_0__inst_mult_5_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_71 (
// Equation(s):
// Xd_0__inst_mult_2_184  = SUM(( !Xd_0__inst_mult_2_6_q  $ (!Xd_0__inst_mult_2_7_q ) ) + ( Xd_0__inst_mult_2_182  ) + ( Xd_0__inst_mult_2_181  ))
// Xd_0__inst_mult_2_185  = CARRY(( !Xd_0__inst_mult_2_6_q  $ (!Xd_0__inst_mult_2_7_q ) ) + ( Xd_0__inst_mult_2_182  ) + ( Xd_0__inst_mult_2_181  ))
// Xd_0__inst_mult_2_186  = SHARE((Xd_0__inst_mult_2_6_q  & Xd_0__inst_mult_2_7_q ))

	.dataa(!Xd_0__inst_mult_2_6_q ),
	.datab(!Xd_0__inst_mult_2_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_181 ),
	.sharein(Xd_0__inst_mult_2_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_184 ),
	.cout(Xd_0__inst_mult_2_185 ),
	.shareout(Xd_0__inst_mult_2_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_67 (
// Equation(s):
// Xd_0__inst_mult_3_180  = SUM(( !Xd_0__inst_mult_3_6_q  $ (!Xd_0__inst_mult_3_7_q ) ) + ( Xd_0__inst_mult_3_178  ) + ( Xd_0__inst_mult_3_177  ))
// Xd_0__inst_mult_3_181  = CARRY(( !Xd_0__inst_mult_3_6_q  $ (!Xd_0__inst_mult_3_7_q ) ) + ( Xd_0__inst_mult_3_178  ) + ( Xd_0__inst_mult_3_177  ))
// Xd_0__inst_mult_3_182  = SHARE((Xd_0__inst_mult_3_6_q  & Xd_0__inst_mult_3_7_q ))

	.dataa(!Xd_0__inst_mult_3_6_q ),
	.datab(!Xd_0__inst_mult_3_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_177 ),
	.sharein(Xd_0__inst_mult_3_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_180 ),
	.cout(Xd_0__inst_mult_3_181 ),
	.shareout(Xd_0__inst_mult_3_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_71 (
// Equation(s):
// Xd_0__inst_mult_0_184  = SUM(( !Xd_0__inst_mult_0_6_q  $ (!Xd_0__inst_mult_0_7_q ) ) + ( Xd_0__inst_mult_0_182  ) + ( Xd_0__inst_mult_0_181  ))
// Xd_0__inst_mult_0_185  = CARRY(( !Xd_0__inst_mult_0_6_q  $ (!Xd_0__inst_mult_0_7_q ) ) + ( Xd_0__inst_mult_0_182  ) + ( Xd_0__inst_mult_0_181  ))
// Xd_0__inst_mult_0_186  = SHARE((Xd_0__inst_mult_0_6_q  & Xd_0__inst_mult_0_7_q ))

	.dataa(!Xd_0__inst_mult_0_6_q ),
	.datab(!Xd_0__inst_mult_0_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_181 ),
	.sharein(Xd_0__inst_mult_0_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_184 ),
	.cout(Xd_0__inst_mult_0_185 ),
	.shareout(Xd_0__inst_mult_0_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_71 (
// Equation(s):
// Xd_0__inst_mult_1_184  = SUM(( !Xd_0__inst_mult_1_6_q  $ (!Xd_0__inst_mult_1_7_q ) ) + ( Xd_0__inst_mult_1_182  ) + ( Xd_0__inst_mult_1_181  ))
// Xd_0__inst_mult_1_185  = CARRY(( !Xd_0__inst_mult_1_6_q  $ (!Xd_0__inst_mult_1_7_q ) ) + ( Xd_0__inst_mult_1_182  ) + ( Xd_0__inst_mult_1_181  ))
// Xd_0__inst_mult_1_186  = SHARE((Xd_0__inst_mult_1_6_q  & Xd_0__inst_mult_1_7_q ))

	.dataa(!Xd_0__inst_mult_1_6_q ),
	.datab(!Xd_0__inst_mult_1_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_181 ),
	.sharein(Xd_0__inst_mult_1_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_184 ),
	.cout(Xd_0__inst_mult_1_185 ),
	.shareout(Xd_0__inst_mult_1_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_74 (
// Equation(s):
// Xd_0__inst_mult_12_208  = SUM(( !Xd_0__inst_mult_12_8_q  $ (!Xd_0__inst_mult_12_9_q ) ) + ( Xd_0__inst_mult_12_206  ) + ( Xd_0__inst_mult_12_205  ))
// Xd_0__inst_mult_12_209  = CARRY(( !Xd_0__inst_mult_12_8_q  $ (!Xd_0__inst_mult_12_9_q ) ) + ( Xd_0__inst_mult_12_206  ) + ( Xd_0__inst_mult_12_205  ))
// Xd_0__inst_mult_12_210  = SHARE((Xd_0__inst_mult_12_8_q  & Xd_0__inst_mult_12_9_q ))

	.dataa(!Xd_0__inst_mult_12_8_q ),
	.datab(!Xd_0__inst_mult_12_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_205 ),
	.sharein(Xd_0__inst_mult_12_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_208 ),
	.cout(Xd_0__inst_mult_12_209 ),
	.shareout(Xd_0__inst_mult_12_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_74 (
// Equation(s):
// Xd_0__inst_mult_13_196  = SUM(( !Xd_0__inst_mult_13_8_q  $ (!Xd_0__inst_mult_13_9_q ) ) + ( Xd_0__inst_mult_13_194  ) + ( Xd_0__inst_mult_13_193  ))
// Xd_0__inst_mult_13_197  = CARRY(( !Xd_0__inst_mult_13_8_q  $ (!Xd_0__inst_mult_13_9_q ) ) + ( Xd_0__inst_mult_13_194  ) + ( Xd_0__inst_mult_13_193  ))
// Xd_0__inst_mult_13_198  = SHARE((Xd_0__inst_mult_13_8_q  & Xd_0__inst_mult_13_9_q ))

	.dataa(!Xd_0__inst_mult_13_8_q ),
	.datab(!Xd_0__inst_mult_13_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_193 ),
	.sharein(Xd_0__inst_mult_13_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_196 ),
	.cout(Xd_0__inst_mult_13_197 ),
	.shareout(Xd_0__inst_mult_13_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_78 (
// Equation(s):
// Xd_0__inst_mult_14_212  = SUM(( !Xd_0__inst_mult_14_8_q  $ (!Xd_0__inst_mult_14_9_q ) ) + ( Xd_0__inst_mult_14_210  ) + ( Xd_0__inst_mult_14_209  ))
// Xd_0__inst_mult_14_213  = CARRY(( !Xd_0__inst_mult_14_8_q  $ (!Xd_0__inst_mult_14_9_q ) ) + ( Xd_0__inst_mult_14_210  ) + ( Xd_0__inst_mult_14_209  ))
// Xd_0__inst_mult_14_214  = SHARE((Xd_0__inst_mult_14_8_q  & Xd_0__inst_mult_14_9_q ))

	.dataa(!Xd_0__inst_mult_14_8_q ),
	.datab(!Xd_0__inst_mult_14_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_209 ),
	.sharein(Xd_0__inst_mult_14_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_212 ),
	.cout(Xd_0__inst_mult_14_213 ),
	.shareout(Xd_0__inst_mult_14_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_78 (
// Equation(s):
// Xd_0__inst_mult_15_212  = SUM(( !Xd_0__inst_mult_15_8_q  $ (!Xd_0__inst_mult_15_9_q ) ) + ( Xd_0__inst_mult_15_210  ) + ( Xd_0__inst_mult_15_209  ))
// Xd_0__inst_mult_15_213  = CARRY(( !Xd_0__inst_mult_15_8_q  $ (!Xd_0__inst_mult_15_9_q ) ) + ( Xd_0__inst_mult_15_210  ) + ( Xd_0__inst_mult_15_209  ))
// Xd_0__inst_mult_15_214  = SHARE((Xd_0__inst_mult_15_8_q  & Xd_0__inst_mult_15_9_q ))

	.dataa(!Xd_0__inst_mult_15_8_q ),
	.datab(!Xd_0__inst_mult_15_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_209 ),
	.sharein(Xd_0__inst_mult_15_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_212 ),
	.cout(Xd_0__inst_mult_15_213 ),
	.shareout(Xd_0__inst_mult_15_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_70 (
// Equation(s):
// Xd_0__inst_mult_10_192  = SUM(( !Xd_0__inst_mult_10_8_q  $ (!Xd_0__inst_mult_10_9_q ) ) + ( Xd_0__inst_mult_10_190  ) + ( Xd_0__inst_mult_10_189  ))
// Xd_0__inst_mult_10_193  = CARRY(( !Xd_0__inst_mult_10_8_q  $ (!Xd_0__inst_mult_10_9_q ) ) + ( Xd_0__inst_mult_10_190  ) + ( Xd_0__inst_mult_10_189  ))
// Xd_0__inst_mult_10_194  = SHARE((Xd_0__inst_mult_10_8_q  & Xd_0__inst_mult_10_9_q ))

	.dataa(!Xd_0__inst_mult_10_8_q ),
	.datab(!Xd_0__inst_mult_10_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_189 ),
	.sharein(Xd_0__inst_mult_10_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_192 ),
	.cout(Xd_0__inst_mult_10_193 ),
	.shareout(Xd_0__inst_mult_10_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_74 (
// Equation(s):
// Xd_0__inst_mult_11_196  = SUM(( !Xd_0__inst_mult_11_8_q  $ (!Xd_0__inst_mult_11_9_q ) ) + ( Xd_0__inst_mult_11_194  ) + ( Xd_0__inst_mult_11_193  ))
// Xd_0__inst_mult_11_197  = CARRY(( !Xd_0__inst_mult_11_8_q  $ (!Xd_0__inst_mult_11_9_q ) ) + ( Xd_0__inst_mult_11_194  ) + ( Xd_0__inst_mult_11_193  ))
// Xd_0__inst_mult_11_198  = SHARE((Xd_0__inst_mult_11_8_q  & Xd_0__inst_mult_11_9_q ))

	.dataa(!Xd_0__inst_mult_11_8_q ),
	.datab(!Xd_0__inst_mult_11_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_193 ),
	.sharein(Xd_0__inst_mult_11_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_196 ),
	.cout(Xd_0__inst_mult_11_197 ),
	.shareout(Xd_0__inst_mult_11_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_74 (
// Equation(s):
// Xd_0__inst_mult_8_196  = SUM(( !Xd_0__inst_mult_8_8_q  $ (!Xd_0__inst_mult_8_9_q ) ) + ( Xd_0__inst_mult_8_194  ) + ( Xd_0__inst_mult_8_193  ))
// Xd_0__inst_mult_8_197  = CARRY(( !Xd_0__inst_mult_8_8_q  $ (!Xd_0__inst_mult_8_9_q ) ) + ( Xd_0__inst_mult_8_194  ) + ( Xd_0__inst_mult_8_193  ))
// Xd_0__inst_mult_8_198  = SHARE((Xd_0__inst_mult_8_8_q  & Xd_0__inst_mult_8_9_q ))

	.dataa(!Xd_0__inst_mult_8_8_q ),
	.datab(!Xd_0__inst_mult_8_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_193 ),
	.sharein(Xd_0__inst_mult_8_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_196 ),
	.cout(Xd_0__inst_mult_8_197 ),
	.shareout(Xd_0__inst_mult_8_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_70 (
// Equation(s):
// Xd_0__inst_mult_9_192  = SUM(( !Xd_0__inst_mult_9_8_q  $ (!Xd_0__inst_mult_9_9_q ) ) + ( Xd_0__inst_mult_9_190  ) + ( Xd_0__inst_mult_9_189  ))
// Xd_0__inst_mult_9_193  = CARRY(( !Xd_0__inst_mult_9_8_q  $ (!Xd_0__inst_mult_9_9_q ) ) + ( Xd_0__inst_mult_9_190  ) + ( Xd_0__inst_mult_9_189  ))
// Xd_0__inst_mult_9_194  = SHARE((Xd_0__inst_mult_9_8_q  & Xd_0__inst_mult_9_9_q ))

	.dataa(!Xd_0__inst_mult_9_8_q ),
	.datab(!Xd_0__inst_mult_9_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_189 ),
	.sharein(Xd_0__inst_mult_9_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_192 ),
	.cout(Xd_0__inst_mult_9_193 ),
	.shareout(Xd_0__inst_mult_9_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_70 (
// Equation(s):
// Xd_0__inst_mult_6_192  = SUM(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q ) ) + ( Xd_0__inst_mult_6_190  ) + ( Xd_0__inst_mult_6_189  ))
// Xd_0__inst_mult_6_193  = CARRY(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q ) ) + ( Xd_0__inst_mult_6_190  ) + ( Xd_0__inst_mult_6_189  ))
// Xd_0__inst_mult_6_194  = SHARE((Xd_0__inst_mult_6_8_q  & Xd_0__inst_mult_6_9_q ))

	.dataa(!Xd_0__inst_mult_6_8_q ),
	.datab(!Xd_0__inst_mult_6_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_189 ),
	.sharein(Xd_0__inst_mult_6_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_192 ),
	.cout(Xd_0__inst_mult_6_193 ),
	.shareout(Xd_0__inst_mult_6_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_68 (
// Equation(s):
// Xd_0__inst_mult_7_184  = SUM(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q ) ) + ( Xd_0__inst_mult_7_182  ) + ( Xd_0__inst_mult_7_181  ))
// Xd_0__inst_mult_7_185  = CARRY(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q ) ) + ( Xd_0__inst_mult_7_182  ) + ( Xd_0__inst_mult_7_181  ))
// Xd_0__inst_mult_7_186  = SHARE((Xd_0__inst_mult_7_8_q  & Xd_0__inst_mult_7_9_q ))

	.dataa(!Xd_0__inst_mult_7_8_q ),
	.datab(!Xd_0__inst_mult_7_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_181 ),
	.sharein(Xd_0__inst_mult_7_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_184 ),
	.cout(Xd_0__inst_mult_7_185 ),
	.shareout(Xd_0__inst_mult_7_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_78 (
// Equation(s):
// Xd_0__inst_mult_4_212  = SUM(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q ) ) + ( Xd_0__inst_mult_4_210  ) + ( Xd_0__inst_mult_4_209  ))
// Xd_0__inst_mult_4_213  = CARRY(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q ) ) + ( Xd_0__inst_mult_4_210  ) + ( Xd_0__inst_mult_4_209  ))
// Xd_0__inst_mult_4_214  = SHARE((Xd_0__inst_mult_4_8_q  & Xd_0__inst_mult_4_9_q ))

	.dataa(!Xd_0__inst_mult_4_8_q ),
	.datab(!Xd_0__inst_mult_4_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_209 ),
	.sharein(Xd_0__inst_mult_4_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_212 ),
	.cout(Xd_0__inst_mult_4_213 ),
	.shareout(Xd_0__inst_mult_4_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_68 (
// Equation(s):
// Xd_0__inst_mult_5_184  = SUM(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q ) ) + ( Xd_0__inst_mult_5_182  ) + ( Xd_0__inst_mult_5_181  ))
// Xd_0__inst_mult_5_185  = CARRY(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q ) ) + ( Xd_0__inst_mult_5_182  ) + ( Xd_0__inst_mult_5_181  ))
// Xd_0__inst_mult_5_186  = SHARE((Xd_0__inst_mult_5_8_q  & Xd_0__inst_mult_5_9_q ))

	.dataa(!Xd_0__inst_mult_5_8_q ),
	.datab(!Xd_0__inst_mult_5_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_181 ),
	.sharein(Xd_0__inst_mult_5_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_184 ),
	.cout(Xd_0__inst_mult_5_185 ),
	.shareout(Xd_0__inst_mult_5_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_72 (
// Equation(s):
// Xd_0__inst_mult_2_188  = SUM(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q ) ) + ( Xd_0__inst_mult_2_186  ) + ( Xd_0__inst_mult_2_185  ))
// Xd_0__inst_mult_2_189  = CARRY(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q ) ) + ( Xd_0__inst_mult_2_186  ) + ( Xd_0__inst_mult_2_185  ))
// Xd_0__inst_mult_2_190  = SHARE((Xd_0__inst_mult_2_8_q  & Xd_0__inst_mult_2_9_q ))

	.dataa(!Xd_0__inst_mult_2_8_q ),
	.datab(!Xd_0__inst_mult_2_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_185 ),
	.sharein(Xd_0__inst_mult_2_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_188 ),
	.cout(Xd_0__inst_mult_2_189 ),
	.shareout(Xd_0__inst_mult_2_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_68 (
// Equation(s):
// Xd_0__inst_mult_3_184  = SUM(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q ) ) + ( Xd_0__inst_mult_3_182  ) + ( Xd_0__inst_mult_3_181  ))
// Xd_0__inst_mult_3_185  = CARRY(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q ) ) + ( Xd_0__inst_mult_3_182  ) + ( Xd_0__inst_mult_3_181  ))
// Xd_0__inst_mult_3_186  = SHARE((Xd_0__inst_mult_3_8_q  & Xd_0__inst_mult_3_9_q ))

	.dataa(!Xd_0__inst_mult_3_8_q ),
	.datab(!Xd_0__inst_mult_3_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_181 ),
	.sharein(Xd_0__inst_mult_3_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_184 ),
	.cout(Xd_0__inst_mult_3_185 ),
	.shareout(Xd_0__inst_mult_3_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_72 (
// Equation(s):
// Xd_0__inst_mult_0_188  = SUM(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q ) ) + ( Xd_0__inst_mult_0_186  ) + ( Xd_0__inst_mult_0_185  ))
// Xd_0__inst_mult_0_189  = CARRY(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q ) ) + ( Xd_0__inst_mult_0_186  ) + ( Xd_0__inst_mult_0_185  ))
// Xd_0__inst_mult_0_190  = SHARE((Xd_0__inst_mult_0_8_q  & Xd_0__inst_mult_0_9_q ))

	.dataa(!Xd_0__inst_mult_0_8_q ),
	.datab(!Xd_0__inst_mult_0_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_185 ),
	.sharein(Xd_0__inst_mult_0_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_188 ),
	.cout(Xd_0__inst_mult_0_189 ),
	.shareout(Xd_0__inst_mult_0_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_72 (
// Equation(s):
// Xd_0__inst_mult_1_188  = SUM(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q ) ) + ( Xd_0__inst_mult_1_186  ) + ( Xd_0__inst_mult_1_185  ))
// Xd_0__inst_mult_1_189  = CARRY(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q ) ) + ( Xd_0__inst_mult_1_186  ) + ( Xd_0__inst_mult_1_185  ))
// Xd_0__inst_mult_1_190  = SHARE((Xd_0__inst_mult_1_8_q  & Xd_0__inst_mult_1_9_q ))

	.dataa(!Xd_0__inst_mult_1_8_q ),
	.datab(!Xd_0__inst_mult_1_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_185 ),
	.sharein(Xd_0__inst_mult_1_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_188 ),
	.cout(Xd_0__inst_mult_1_189 ),
	.shareout(Xd_0__inst_mult_1_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_75 (
// Equation(s):
// Xd_0__inst_mult_12_212  = SUM(( !Xd_0__inst_mult_12_10_q  $ (!Xd_0__inst_mult_12_11_q ) ) + ( Xd_0__inst_mult_12_210  ) + ( Xd_0__inst_mult_12_209  ))
// Xd_0__inst_mult_12_213  = CARRY(( !Xd_0__inst_mult_12_10_q  $ (!Xd_0__inst_mult_12_11_q ) ) + ( Xd_0__inst_mult_12_210  ) + ( Xd_0__inst_mult_12_209  ))
// Xd_0__inst_mult_12_214  = SHARE((Xd_0__inst_mult_12_10_q  & Xd_0__inst_mult_12_11_q ))

	.dataa(!Xd_0__inst_mult_12_10_q ),
	.datab(!Xd_0__inst_mult_12_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_209 ),
	.sharein(Xd_0__inst_mult_12_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_212 ),
	.cout(Xd_0__inst_mult_12_213 ),
	.shareout(Xd_0__inst_mult_12_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_75 (
// Equation(s):
// Xd_0__inst_mult_13_200  = SUM(( !Xd_0__inst_mult_13_10_q  $ (!Xd_0__inst_mult_13_11_q ) ) + ( Xd_0__inst_mult_13_198  ) + ( Xd_0__inst_mult_13_197  ))
// Xd_0__inst_mult_13_201  = CARRY(( !Xd_0__inst_mult_13_10_q  $ (!Xd_0__inst_mult_13_11_q ) ) + ( Xd_0__inst_mult_13_198  ) + ( Xd_0__inst_mult_13_197  ))
// Xd_0__inst_mult_13_202  = SHARE((Xd_0__inst_mult_13_10_q  & Xd_0__inst_mult_13_11_q ))

	.dataa(!Xd_0__inst_mult_13_10_q ),
	.datab(!Xd_0__inst_mult_13_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_197 ),
	.sharein(Xd_0__inst_mult_13_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_200 ),
	.cout(Xd_0__inst_mult_13_201 ),
	.shareout(Xd_0__inst_mult_13_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_79 (
// Equation(s):
// Xd_0__inst_mult_14_216  = SUM(( !Xd_0__inst_mult_14_10_q  $ (!Xd_0__inst_mult_14_11_q ) ) + ( Xd_0__inst_mult_14_214  ) + ( Xd_0__inst_mult_14_213  ))
// Xd_0__inst_mult_14_217  = CARRY(( !Xd_0__inst_mult_14_10_q  $ (!Xd_0__inst_mult_14_11_q ) ) + ( Xd_0__inst_mult_14_214  ) + ( Xd_0__inst_mult_14_213  ))
// Xd_0__inst_mult_14_218  = SHARE((Xd_0__inst_mult_14_10_q  & Xd_0__inst_mult_14_11_q ))

	.dataa(!Xd_0__inst_mult_14_10_q ),
	.datab(!Xd_0__inst_mult_14_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_213 ),
	.sharein(Xd_0__inst_mult_14_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_216 ),
	.cout(Xd_0__inst_mult_14_217 ),
	.shareout(Xd_0__inst_mult_14_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_79 (
// Equation(s):
// Xd_0__inst_mult_15_216  = SUM(( !Xd_0__inst_mult_15_10_q  $ (!Xd_0__inst_mult_15_11_q ) ) + ( Xd_0__inst_mult_15_214  ) + ( Xd_0__inst_mult_15_213  ))
// Xd_0__inst_mult_15_217  = CARRY(( !Xd_0__inst_mult_15_10_q  $ (!Xd_0__inst_mult_15_11_q ) ) + ( Xd_0__inst_mult_15_214  ) + ( Xd_0__inst_mult_15_213  ))
// Xd_0__inst_mult_15_218  = SHARE((Xd_0__inst_mult_15_10_q  & Xd_0__inst_mult_15_11_q ))

	.dataa(!Xd_0__inst_mult_15_10_q ),
	.datab(!Xd_0__inst_mult_15_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_213 ),
	.sharein(Xd_0__inst_mult_15_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_216 ),
	.cout(Xd_0__inst_mult_15_217 ),
	.shareout(Xd_0__inst_mult_15_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_71 (
// Equation(s):
// Xd_0__inst_mult_10_196  = SUM(( !Xd_0__inst_mult_10_10_q  $ (!Xd_0__inst_mult_10_11_q ) ) + ( Xd_0__inst_mult_10_194  ) + ( Xd_0__inst_mult_10_193  ))
// Xd_0__inst_mult_10_197  = CARRY(( !Xd_0__inst_mult_10_10_q  $ (!Xd_0__inst_mult_10_11_q ) ) + ( Xd_0__inst_mult_10_194  ) + ( Xd_0__inst_mult_10_193  ))
// Xd_0__inst_mult_10_198  = SHARE((Xd_0__inst_mult_10_10_q  & Xd_0__inst_mult_10_11_q ))

	.dataa(!Xd_0__inst_mult_10_10_q ),
	.datab(!Xd_0__inst_mult_10_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_193 ),
	.sharein(Xd_0__inst_mult_10_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_196 ),
	.cout(Xd_0__inst_mult_10_197 ),
	.shareout(Xd_0__inst_mult_10_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_75 (
// Equation(s):
// Xd_0__inst_mult_11_200  = SUM(( !Xd_0__inst_mult_11_10_q  $ (!Xd_0__inst_mult_11_11_q ) ) + ( Xd_0__inst_mult_11_198  ) + ( Xd_0__inst_mult_11_197  ))
// Xd_0__inst_mult_11_201  = CARRY(( !Xd_0__inst_mult_11_10_q  $ (!Xd_0__inst_mult_11_11_q ) ) + ( Xd_0__inst_mult_11_198  ) + ( Xd_0__inst_mult_11_197  ))
// Xd_0__inst_mult_11_202  = SHARE((Xd_0__inst_mult_11_10_q  & Xd_0__inst_mult_11_11_q ))

	.dataa(!Xd_0__inst_mult_11_10_q ),
	.datab(!Xd_0__inst_mult_11_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_197 ),
	.sharein(Xd_0__inst_mult_11_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_200 ),
	.cout(Xd_0__inst_mult_11_201 ),
	.shareout(Xd_0__inst_mult_11_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_75 (
// Equation(s):
// Xd_0__inst_mult_8_200  = SUM(( !Xd_0__inst_mult_8_10_q  $ (!Xd_0__inst_mult_8_11_q ) ) + ( Xd_0__inst_mult_8_198  ) + ( Xd_0__inst_mult_8_197  ))
// Xd_0__inst_mult_8_201  = CARRY(( !Xd_0__inst_mult_8_10_q  $ (!Xd_0__inst_mult_8_11_q ) ) + ( Xd_0__inst_mult_8_198  ) + ( Xd_0__inst_mult_8_197  ))
// Xd_0__inst_mult_8_202  = SHARE((Xd_0__inst_mult_8_10_q  & Xd_0__inst_mult_8_11_q ))

	.dataa(!Xd_0__inst_mult_8_10_q ),
	.datab(!Xd_0__inst_mult_8_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_197 ),
	.sharein(Xd_0__inst_mult_8_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_200 ),
	.cout(Xd_0__inst_mult_8_201 ),
	.shareout(Xd_0__inst_mult_8_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_71 (
// Equation(s):
// Xd_0__inst_mult_9_196  = SUM(( !Xd_0__inst_mult_9_10_q  $ (!Xd_0__inst_mult_9_11_q ) ) + ( Xd_0__inst_mult_9_194  ) + ( Xd_0__inst_mult_9_193  ))
// Xd_0__inst_mult_9_197  = CARRY(( !Xd_0__inst_mult_9_10_q  $ (!Xd_0__inst_mult_9_11_q ) ) + ( Xd_0__inst_mult_9_194  ) + ( Xd_0__inst_mult_9_193  ))
// Xd_0__inst_mult_9_198  = SHARE((Xd_0__inst_mult_9_10_q  & Xd_0__inst_mult_9_11_q ))

	.dataa(!Xd_0__inst_mult_9_10_q ),
	.datab(!Xd_0__inst_mult_9_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_193 ),
	.sharein(Xd_0__inst_mult_9_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_196 ),
	.cout(Xd_0__inst_mult_9_197 ),
	.shareout(Xd_0__inst_mult_9_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_71 (
// Equation(s):
// Xd_0__inst_mult_6_196  = SUM(( !Xd_0__inst_mult_6_10_q  $ (!Xd_0__inst_mult_6_11_q ) ) + ( Xd_0__inst_mult_6_194  ) + ( Xd_0__inst_mult_6_193  ))
// Xd_0__inst_mult_6_197  = CARRY(( !Xd_0__inst_mult_6_10_q  $ (!Xd_0__inst_mult_6_11_q ) ) + ( Xd_0__inst_mult_6_194  ) + ( Xd_0__inst_mult_6_193  ))
// Xd_0__inst_mult_6_198  = SHARE((Xd_0__inst_mult_6_10_q  & Xd_0__inst_mult_6_11_q ))

	.dataa(!Xd_0__inst_mult_6_10_q ),
	.datab(!Xd_0__inst_mult_6_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_193 ),
	.sharein(Xd_0__inst_mult_6_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_196 ),
	.cout(Xd_0__inst_mult_6_197 ),
	.shareout(Xd_0__inst_mult_6_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_69 (
// Equation(s):
// Xd_0__inst_mult_7_188  = SUM(( !Xd_0__inst_mult_7_10_q  $ (!Xd_0__inst_mult_7_11_q ) ) + ( Xd_0__inst_mult_7_186  ) + ( Xd_0__inst_mult_7_185  ))
// Xd_0__inst_mult_7_189  = CARRY(( !Xd_0__inst_mult_7_10_q  $ (!Xd_0__inst_mult_7_11_q ) ) + ( Xd_0__inst_mult_7_186  ) + ( Xd_0__inst_mult_7_185  ))
// Xd_0__inst_mult_7_190  = SHARE((Xd_0__inst_mult_7_10_q  & Xd_0__inst_mult_7_11_q ))

	.dataa(!Xd_0__inst_mult_7_10_q ),
	.datab(!Xd_0__inst_mult_7_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_185 ),
	.sharein(Xd_0__inst_mult_7_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_188 ),
	.cout(Xd_0__inst_mult_7_189 ),
	.shareout(Xd_0__inst_mult_7_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_79 (
// Equation(s):
// Xd_0__inst_mult_4_216  = SUM(( !Xd_0__inst_mult_4_10_q  $ (!Xd_0__inst_mult_4_11_q ) ) + ( Xd_0__inst_mult_4_214  ) + ( Xd_0__inst_mult_4_213  ))
// Xd_0__inst_mult_4_217  = CARRY(( !Xd_0__inst_mult_4_10_q  $ (!Xd_0__inst_mult_4_11_q ) ) + ( Xd_0__inst_mult_4_214  ) + ( Xd_0__inst_mult_4_213  ))
// Xd_0__inst_mult_4_218  = SHARE((Xd_0__inst_mult_4_10_q  & Xd_0__inst_mult_4_11_q ))

	.dataa(!Xd_0__inst_mult_4_10_q ),
	.datab(!Xd_0__inst_mult_4_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_213 ),
	.sharein(Xd_0__inst_mult_4_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_216 ),
	.cout(Xd_0__inst_mult_4_217 ),
	.shareout(Xd_0__inst_mult_4_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_69 (
// Equation(s):
// Xd_0__inst_mult_5_188  = SUM(( !Xd_0__inst_mult_5_10_q  $ (!Xd_0__inst_mult_5_11_q ) ) + ( Xd_0__inst_mult_5_186  ) + ( Xd_0__inst_mult_5_185  ))
// Xd_0__inst_mult_5_189  = CARRY(( !Xd_0__inst_mult_5_10_q  $ (!Xd_0__inst_mult_5_11_q ) ) + ( Xd_0__inst_mult_5_186  ) + ( Xd_0__inst_mult_5_185  ))
// Xd_0__inst_mult_5_190  = SHARE((Xd_0__inst_mult_5_10_q  & Xd_0__inst_mult_5_11_q ))

	.dataa(!Xd_0__inst_mult_5_10_q ),
	.datab(!Xd_0__inst_mult_5_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_185 ),
	.sharein(Xd_0__inst_mult_5_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_188 ),
	.cout(Xd_0__inst_mult_5_189 ),
	.shareout(Xd_0__inst_mult_5_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_73 (
// Equation(s):
// Xd_0__inst_mult_2_192  = SUM(( !Xd_0__inst_mult_2_10_q  $ (!Xd_0__inst_mult_2_11_q ) ) + ( Xd_0__inst_mult_2_190  ) + ( Xd_0__inst_mult_2_189  ))
// Xd_0__inst_mult_2_193  = CARRY(( !Xd_0__inst_mult_2_10_q  $ (!Xd_0__inst_mult_2_11_q ) ) + ( Xd_0__inst_mult_2_190  ) + ( Xd_0__inst_mult_2_189  ))
// Xd_0__inst_mult_2_194  = SHARE((Xd_0__inst_mult_2_10_q  & Xd_0__inst_mult_2_11_q ))

	.dataa(!Xd_0__inst_mult_2_10_q ),
	.datab(!Xd_0__inst_mult_2_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_189 ),
	.sharein(Xd_0__inst_mult_2_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_192 ),
	.cout(Xd_0__inst_mult_2_193 ),
	.shareout(Xd_0__inst_mult_2_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_69 (
// Equation(s):
// Xd_0__inst_mult_3_188  = SUM(( !Xd_0__inst_mult_3_10_q  $ (!Xd_0__inst_mult_3_11_q ) ) + ( Xd_0__inst_mult_3_186  ) + ( Xd_0__inst_mult_3_185  ))
// Xd_0__inst_mult_3_189  = CARRY(( !Xd_0__inst_mult_3_10_q  $ (!Xd_0__inst_mult_3_11_q ) ) + ( Xd_0__inst_mult_3_186  ) + ( Xd_0__inst_mult_3_185  ))
// Xd_0__inst_mult_3_190  = SHARE((Xd_0__inst_mult_3_10_q  & Xd_0__inst_mult_3_11_q ))

	.dataa(!Xd_0__inst_mult_3_10_q ),
	.datab(!Xd_0__inst_mult_3_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_185 ),
	.sharein(Xd_0__inst_mult_3_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_188 ),
	.cout(Xd_0__inst_mult_3_189 ),
	.shareout(Xd_0__inst_mult_3_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_73 (
// Equation(s):
// Xd_0__inst_mult_0_192  = SUM(( !Xd_0__inst_mult_0_10_q  $ (!Xd_0__inst_mult_0_11_q ) ) + ( Xd_0__inst_mult_0_190  ) + ( Xd_0__inst_mult_0_189  ))
// Xd_0__inst_mult_0_193  = CARRY(( !Xd_0__inst_mult_0_10_q  $ (!Xd_0__inst_mult_0_11_q ) ) + ( Xd_0__inst_mult_0_190  ) + ( Xd_0__inst_mult_0_189  ))
// Xd_0__inst_mult_0_194  = SHARE((Xd_0__inst_mult_0_10_q  & Xd_0__inst_mult_0_11_q ))

	.dataa(!Xd_0__inst_mult_0_10_q ),
	.datab(!Xd_0__inst_mult_0_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_189 ),
	.sharein(Xd_0__inst_mult_0_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_192 ),
	.cout(Xd_0__inst_mult_0_193 ),
	.shareout(Xd_0__inst_mult_0_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_73 (
// Equation(s):
// Xd_0__inst_mult_1_192  = SUM(( !Xd_0__inst_mult_1_10_q  $ (!Xd_0__inst_mult_1_11_q ) ) + ( Xd_0__inst_mult_1_190  ) + ( Xd_0__inst_mult_1_189  ))
// Xd_0__inst_mult_1_193  = CARRY(( !Xd_0__inst_mult_1_10_q  $ (!Xd_0__inst_mult_1_11_q ) ) + ( Xd_0__inst_mult_1_190  ) + ( Xd_0__inst_mult_1_189  ))
// Xd_0__inst_mult_1_194  = SHARE((Xd_0__inst_mult_1_10_q  & Xd_0__inst_mult_1_11_q ))

	.dataa(!Xd_0__inst_mult_1_10_q ),
	.datab(!Xd_0__inst_mult_1_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_189 ),
	.sharein(Xd_0__inst_mult_1_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_192 ),
	.cout(Xd_0__inst_mult_1_193 ),
	.shareout(Xd_0__inst_mult_1_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_76 (
// Equation(s):
// Xd_0__inst_mult_12_216  = SUM(( !Xd_0__inst_mult_12_12_q  $ (!Xd_0__inst_mult_12_13_q ) ) + ( Xd_0__inst_mult_12_214  ) + ( Xd_0__inst_mult_12_213  ))
// Xd_0__inst_mult_12_217  = CARRY(( !Xd_0__inst_mult_12_12_q  $ (!Xd_0__inst_mult_12_13_q ) ) + ( Xd_0__inst_mult_12_214  ) + ( Xd_0__inst_mult_12_213  ))
// Xd_0__inst_mult_12_218  = SHARE((Xd_0__inst_mult_12_12_q  & Xd_0__inst_mult_12_13_q ))

	.dataa(!Xd_0__inst_mult_12_12_q ),
	.datab(!Xd_0__inst_mult_12_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_213 ),
	.sharein(Xd_0__inst_mult_12_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_216 ),
	.cout(Xd_0__inst_mult_12_217 ),
	.shareout(Xd_0__inst_mult_12_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_76 (
// Equation(s):
// Xd_0__inst_mult_13_204  = SUM(( !Xd_0__inst_mult_13_12_q  $ (!Xd_0__inst_mult_13_13_q ) ) + ( Xd_0__inst_mult_13_202  ) + ( Xd_0__inst_mult_13_201  ))
// Xd_0__inst_mult_13_205  = CARRY(( !Xd_0__inst_mult_13_12_q  $ (!Xd_0__inst_mult_13_13_q ) ) + ( Xd_0__inst_mult_13_202  ) + ( Xd_0__inst_mult_13_201  ))
// Xd_0__inst_mult_13_206  = SHARE((Xd_0__inst_mult_13_12_q  & Xd_0__inst_mult_13_13_q ))

	.dataa(!Xd_0__inst_mult_13_12_q ),
	.datab(!Xd_0__inst_mult_13_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_201 ),
	.sharein(Xd_0__inst_mult_13_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_204 ),
	.cout(Xd_0__inst_mult_13_205 ),
	.shareout(Xd_0__inst_mult_13_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_80 (
// Equation(s):
// Xd_0__inst_mult_14_220  = SUM(( !Xd_0__inst_mult_14_12_q  $ (!Xd_0__inst_mult_14_13_q ) ) + ( Xd_0__inst_mult_14_218  ) + ( Xd_0__inst_mult_14_217  ))
// Xd_0__inst_mult_14_221  = CARRY(( !Xd_0__inst_mult_14_12_q  $ (!Xd_0__inst_mult_14_13_q ) ) + ( Xd_0__inst_mult_14_218  ) + ( Xd_0__inst_mult_14_217  ))
// Xd_0__inst_mult_14_222  = SHARE((Xd_0__inst_mult_14_12_q  & Xd_0__inst_mult_14_13_q ))

	.dataa(!Xd_0__inst_mult_14_12_q ),
	.datab(!Xd_0__inst_mult_14_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_217 ),
	.sharein(Xd_0__inst_mult_14_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_220 ),
	.cout(Xd_0__inst_mult_14_221 ),
	.shareout(Xd_0__inst_mult_14_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_80 (
// Equation(s):
// Xd_0__inst_mult_15_220  = SUM(( !Xd_0__inst_mult_15_12_q  $ (!Xd_0__inst_mult_15_13_q ) ) + ( Xd_0__inst_mult_15_218  ) + ( Xd_0__inst_mult_15_217  ))
// Xd_0__inst_mult_15_221  = CARRY(( !Xd_0__inst_mult_15_12_q  $ (!Xd_0__inst_mult_15_13_q ) ) + ( Xd_0__inst_mult_15_218  ) + ( Xd_0__inst_mult_15_217  ))
// Xd_0__inst_mult_15_222  = SHARE((Xd_0__inst_mult_15_12_q  & Xd_0__inst_mult_15_13_q ))

	.dataa(!Xd_0__inst_mult_15_12_q ),
	.datab(!Xd_0__inst_mult_15_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_217 ),
	.sharein(Xd_0__inst_mult_15_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_220 ),
	.cout(Xd_0__inst_mult_15_221 ),
	.shareout(Xd_0__inst_mult_15_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_72 (
// Equation(s):
// Xd_0__inst_mult_10_200  = SUM(( !Xd_0__inst_mult_10_12_q  $ (!Xd_0__inst_mult_10_13_q ) ) + ( Xd_0__inst_mult_10_198  ) + ( Xd_0__inst_mult_10_197  ))
// Xd_0__inst_mult_10_201  = CARRY(( !Xd_0__inst_mult_10_12_q  $ (!Xd_0__inst_mult_10_13_q ) ) + ( Xd_0__inst_mult_10_198  ) + ( Xd_0__inst_mult_10_197  ))
// Xd_0__inst_mult_10_202  = SHARE((Xd_0__inst_mult_10_12_q  & Xd_0__inst_mult_10_13_q ))

	.dataa(!Xd_0__inst_mult_10_12_q ),
	.datab(!Xd_0__inst_mult_10_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_197 ),
	.sharein(Xd_0__inst_mult_10_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_200 ),
	.cout(Xd_0__inst_mult_10_201 ),
	.shareout(Xd_0__inst_mult_10_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_76 (
// Equation(s):
// Xd_0__inst_mult_11_204  = SUM(( !Xd_0__inst_mult_11_12_q  $ (!Xd_0__inst_mult_11_13_q ) ) + ( Xd_0__inst_mult_11_202  ) + ( Xd_0__inst_mult_11_201  ))
// Xd_0__inst_mult_11_205  = CARRY(( !Xd_0__inst_mult_11_12_q  $ (!Xd_0__inst_mult_11_13_q ) ) + ( Xd_0__inst_mult_11_202  ) + ( Xd_0__inst_mult_11_201  ))
// Xd_0__inst_mult_11_206  = SHARE((Xd_0__inst_mult_11_12_q  & Xd_0__inst_mult_11_13_q ))

	.dataa(!Xd_0__inst_mult_11_12_q ),
	.datab(!Xd_0__inst_mult_11_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_201 ),
	.sharein(Xd_0__inst_mult_11_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_204 ),
	.cout(Xd_0__inst_mult_11_205 ),
	.shareout(Xd_0__inst_mult_11_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_76 (
// Equation(s):
// Xd_0__inst_mult_8_204  = SUM(( !Xd_0__inst_mult_8_12_q  $ (!Xd_0__inst_mult_8_13_q ) ) + ( Xd_0__inst_mult_8_202  ) + ( Xd_0__inst_mult_8_201  ))
// Xd_0__inst_mult_8_205  = CARRY(( !Xd_0__inst_mult_8_12_q  $ (!Xd_0__inst_mult_8_13_q ) ) + ( Xd_0__inst_mult_8_202  ) + ( Xd_0__inst_mult_8_201  ))
// Xd_0__inst_mult_8_206  = SHARE((Xd_0__inst_mult_8_12_q  & Xd_0__inst_mult_8_13_q ))

	.dataa(!Xd_0__inst_mult_8_12_q ),
	.datab(!Xd_0__inst_mult_8_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_201 ),
	.sharein(Xd_0__inst_mult_8_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_204 ),
	.cout(Xd_0__inst_mult_8_205 ),
	.shareout(Xd_0__inst_mult_8_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_72 (
// Equation(s):
// Xd_0__inst_mult_9_200  = SUM(( !Xd_0__inst_mult_9_12_q  $ (!Xd_0__inst_mult_9_13_q ) ) + ( Xd_0__inst_mult_9_198  ) + ( Xd_0__inst_mult_9_197  ))
// Xd_0__inst_mult_9_201  = CARRY(( !Xd_0__inst_mult_9_12_q  $ (!Xd_0__inst_mult_9_13_q ) ) + ( Xd_0__inst_mult_9_198  ) + ( Xd_0__inst_mult_9_197  ))
// Xd_0__inst_mult_9_202  = SHARE((Xd_0__inst_mult_9_12_q  & Xd_0__inst_mult_9_13_q ))

	.dataa(!Xd_0__inst_mult_9_12_q ),
	.datab(!Xd_0__inst_mult_9_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_197 ),
	.sharein(Xd_0__inst_mult_9_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_200 ),
	.cout(Xd_0__inst_mult_9_201 ),
	.shareout(Xd_0__inst_mult_9_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_72 (
// Equation(s):
// Xd_0__inst_mult_6_200  = SUM(( !Xd_0__inst_mult_6_12_q  $ (!Xd_0__inst_mult_6_13_q ) ) + ( Xd_0__inst_mult_6_198  ) + ( Xd_0__inst_mult_6_197  ))
// Xd_0__inst_mult_6_201  = CARRY(( !Xd_0__inst_mult_6_12_q  $ (!Xd_0__inst_mult_6_13_q ) ) + ( Xd_0__inst_mult_6_198  ) + ( Xd_0__inst_mult_6_197  ))
// Xd_0__inst_mult_6_202  = SHARE((Xd_0__inst_mult_6_12_q  & Xd_0__inst_mult_6_13_q ))

	.dataa(!Xd_0__inst_mult_6_12_q ),
	.datab(!Xd_0__inst_mult_6_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_197 ),
	.sharein(Xd_0__inst_mult_6_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_200 ),
	.cout(Xd_0__inst_mult_6_201 ),
	.shareout(Xd_0__inst_mult_6_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_70 (
// Equation(s):
// Xd_0__inst_mult_7_192  = SUM(( !Xd_0__inst_mult_7_12_q  $ (!Xd_0__inst_mult_7_13_q ) ) + ( Xd_0__inst_mult_7_190  ) + ( Xd_0__inst_mult_7_189  ))
// Xd_0__inst_mult_7_193  = CARRY(( !Xd_0__inst_mult_7_12_q  $ (!Xd_0__inst_mult_7_13_q ) ) + ( Xd_0__inst_mult_7_190  ) + ( Xd_0__inst_mult_7_189  ))
// Xd_0__inst_mult_7_194  = SHARE((Xd_0__inst_mult_7_12_q  & Xd_0__inst_mult_7_13_q ))

	.dataa(!Xd_0__inst_mult_7_12_q ),
	.datab(!Xd_0__inst_mult_7_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_189 ),
	.sharein(Xd_0__inst_mult_7_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_192 ),
	.cout(Xd_0__inst_mult_7_193 ),
	.shareout(Xd_0__inst_mult_7_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_80 (
// Equation(s):
// Xd_0__inst_mult_4_220  = SUM(( !Xd_0__inst_mult_4_12_q  $ (!Xd_0__inst_mult_4_13_q ) ) + ( Xd_0__inst_mult_4_218  ) + ( Xd_0__inst_mult_4_217  ))
// Xd_0__inst_mult_4_221  = CARRY(( !Xd_0__inst_mult_4_12_q  $ (!Xd_0__inst_mult_4_13_q ) ) + ( Xd_0__inst_mult_4_218  ) + ( Xd_0__inst_mult_4_217  ))
// Xd_0__inst_mult_4_222  = SHARE((Xd_0__inst_mult_4_12_q  & Xd_0__inst_mult_4_13_q ))

	.dataa(!Xd_0__inst_mult_4_12_q ),
	.datab(!Xd_0__inst_mult_4_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_217 ),
	.sharein(Xd_0__inst_mult_4_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_220 ),
	.cout(Xd_0__inst_mult_4_221 ),
	.shareout(Xd_0__inst_mult_4_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_70 (
// Equation(s):
// Xd_0__inst_mult_5_192  = SUM(( !Xd_0__inst_mult_5_12_q  $ (!Xd_0__inst_mult_5_13_q ) ) + ( Xd_0__inst_mult_5_190  ) + ( Xd_0__inst_mult_5_189  ))
// Xd_0__inst_mult_5_193  = CARRY(( !Xd_0__inst_mult_5_12_q  $ (!Xd_0__inst_mult_5_13_q ) ) + ( Xd_0__inst_mult_5_190  ) + ( Xd_0__inst_mult_5_189  ))
// Xd_0__inst_mult_5_194  = SHARE((Xd_0__inst_mult_5_12_q  & Xd_0__inst_mult_5_13_q ))

	.dataa(!Xd_0__inst_mult_5_12_q ),
	.datab(!Xd_0__inst_mult_5_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_189 ),
	.sharein(Xd_0__inst_mult_5_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_192 ),
	.cout(Xd_0__inst_mult_5_193 ),
	.shareout(Xd_0__inst_mult_5_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_74 (
// Equation(s):
// Xd_0__inst_mult_2_196  = SUM(( !Xd_0__inst_mult_2_12_q  $ (!Xd_0__inst_mult_2_13_q ) ) + ( Xd_0__inst_mult_2_194  ) + ( Xd_0__inst_mult_2_193  ))
// Xd_0__inst_mult_2_197  = CARRY(( !Xd_0__inst_mult_2_12_q  $ (!Xd_0__inst_mult_2_13_q ) ) + ( Xd_0__inst_mult_2_194  ) + ( Xd_0__inst_mult_2_193  ))
// Xd_0__inst_mult_2_198  = SHARE((Xd_0__inst_mult_2_12_q  & Xd_0__inst_mult_2_13_q ))

	.dataa(!Xd_0__inst_mult_2_12_q ),
	.datab(!Xd_0__inst_mult_2_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_193 ),
	.sharein(Xd_0__inst_mult_2_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_196 ),
	.cout(Xd_0__inst_mult_2_197 ),
	.shareout(Xd_0__inst_mult_2_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_70 (
// Equation(s):
// Xd_0__inst_mult_3_192  = SUM(( !Xd_0__inst_mult_3_12_q  $ (!Xd_0__inst_mult_3_13_q ) ) + ( Xd_0__inst_mult_3_190  ) + ( Xd_0__inst_mult_3_189  ))
// Xd_0__inst_mult_3_193  = CARRY(( !Xd_0__inst_mult_3_12_q  $ (!Xd_0__inst_mult_3_13_q ) ) + ( Xd_0__inst_mult_3_190  ) + ( Xd_0__inst_mult_3_189  ))
// Xd_0__inst_mult_3_194  = SHARE((Xd_0__inst_mult_3_12_q  & Xd_0__inst_mult_3_13_q ))

	.dataa(!Xd_0__inst_mult_3_12_q ),
	.datab(!Xd_0__inst_mult_3_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_189 ),
	.sharein(Xd_0__inst_mult_3_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_192 ),
	.cout(Xd_0__inst_mult_3_193 ),
	.shareout(Xd_0__inst_mult_3_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_74 (
// Equation(s):
// Xd_0__inst_mult_0_196  = SUM(( !Xd_0__inst_mult_0_12_q  $ (!Xd_0__inst_mult_0_13_q ) ) + ( Xd_0__inst_mult_0_194  ) + ( Xd_0__inst_mult_0_193  ))
// Xd_0__inst_mult_0_197  = CARRY(( !Xd_0__inst_mult_0_12_q  $ (!Xd_0__inst_mult_0_13_q ) ) + ( Xd_0__inst_mult_0_194  ) + ( Xd_0__inst_mult_0_193  ))
// Xd_0__inst_mult_0_198  = SHARE((Xd_0__inst_mult_0_12_q  & Xd_0__inst_mult_0_13_q ))

	.dataa(!Xd_0__inst_mult_0_12_q ),
	.datab(!Xd_0__inst_mult_0_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_193 ),
	.sharein(Xd_0__inst_mult_0_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_196 ),
	.cout(Xd_0__inst_mult_0_197 ),
	.shareout(Xd_0__inst_mult_0_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_74 (
// Equation(s):
// Xd_0__inst_mult_1_196  = SUM(( !Xd_0__inst_mult_1_12_q  $ (!Xd_0__inst_mult_1_13_q ) ) + ( Xd_0__inst_mult_1_194  ) + ( Xd_0__inst_mult_1_193  ))
// Xd_0__inst_mult_1_197  = CARRY(( !Xd_0__inst_mult_1_12_q  $ (!Xd_0__inst_mult_1_13_q ) ) + ( Xd_0__inst_mult_1_194  ) + ( Xd_0__inst_mult_1_193  ))
// Xd_0__inst_mult_1_198  = SHARE((Xd_0__inst_mult_1_12_q  & Xd_0__inst_mult_1_13_q ))

	.dataa(!Xd_0__inst_mult_1_12_q ),
	.datab(!Xd_0__inst_mult_1_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_193 ),
	.sharein(Xd_0__inst_mult_1_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_196 ),
	.cout(Xd_0__inst_mult_1_197 ),
	.shareout(Xd_0__inst_mult_1_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_77 (
// Equation(s):
// Xd_0__inst_mult_12_220  = SUM(( !Xd_0__inst_mult_12_14_q  $ (!Xd_0__inst_mult_12_15_q ) ) + ( Xd_0__inst_mult_12_218  ) + ( Xd_0__inst_mult_12_217  ))
// Xd_0__inst_mult_12_221  = CARRY(( !Xd_0__inst_mult_12_14_q  $ (!Xd_0__inst_mult_12_15_q ) ) + ( Xd_0__inst_mult_12_218  ) + ( Xd_0__inst_mult_12_217  ))
// Xd_0__inst_mult_12_222  = SHARE((Xd_0__inst_mult_12_14_q  & Xd_0__inst_mult_12_15_q ))

	.dataa(!Xd_0__inst_mult_12_14_q ),
	.datab(!Xd_0__inst_mult_12_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_217 ),
	.sharein(Xd_0__inst_mult_12_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_220 ),
	.cout(Xd_0__inst_mult_12_221 ),
	.shareout(Xd_0__inst_mult_12_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_77 (
// Equation(s):
// Xd_0__inst_mult_13_208  = SUM(( !Xd_0__inst_mult_13_14_q  $ (!Xd_0__inst_mult_13_15_q ) ) + ( Xd_0__inst_mult_13_206  ) + ( Xd_0__inst_mult_13_205  ))
// Xd_0__inst_mult_13_209  = CARRY(( !Xd_0__inst_mult_13_14_q  $ (!Xd_0__inst_mult_13_15_q ) ) + ( Xd_0__inst_mult_13_206  ) + ( Xd_0__inst_mult_13_205  ))
// Xd_0__inst_mult_13_210  = SHARE((Xd_0__inst_mult_13_14_q  & Xd_0__inst_mult_13_15_q ))

	.dataa(!Xd_0__inst_mult_13_14_q ),
	.datab(!Xd_0__inst_mult_13_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_205 ),
	.sharein(Xd_0__inst_mult_13_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_208 ),
	.cout(Xd_0__inst_mult_13_209 ),
	.shareout(Xd_0__inst_mult_13_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_81 (
// Equation(s):
// Xd_0__inst_mult_14_224  = SUM(( !Xd_0__inst_mult_14_14_q  $ (!Xd_0__inst_mult_14_15_q ) ) + ( Xd_0__inst_mult_14_222  ) + ( Xd_0__inst_mult_14_221  ))
// Xd_0__inst_mult_14_225  = CARRY(( !Xd_0__inst_mult_14_14_q  $ (!Xd_0__inst_mult_14_15_q ) ) + ( Xd_0__inst_mult_14_222  ) + ( Xd_0__inst_mult_14_221  ))
// Xd_0__inst_mult_14_226  = SHARE((Xd_0__inst_mult_14_14_q  & Xd_0__inst_mult_14_15_q ))

	.dataa(!Xd_0__inst_mult_14_14_q ),
	.datab(!Xd_0__inst_mult_14_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_221 ),
	.sharein(Xd_0__inst_mult_14_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_224 ),
	.cout(Xd_0__inst_mult_14_225 ),
	.shareout(Xd_0__inst_mult_14_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_81 (
// Equation(s):
// Xd_0__inst_mult_15_224  = SUM(( !Xd_0__inst_mult_15_14_q  $ (!Xd_0__inst_mult_15_15_q ) ) + ( Xd_0__inst_mult_15_222  ) + ( Xd_0__inst_mult_15_221  ))
// Xd_0__inst_mult_15_225  = CARRY(( !Xd_0__inst_mult_15_14_q  $ (!Xd_0__inst_mult_15_15_q ) ) + ( Xd_0__inst_mult_15_222  ) + ( Xd_0__inst_mult_15_221  ))
// Xd_0__inst_mult_15_226  = SHARE((Xd_0__inst_mult_15_14_q  & Xd_0__inst_mult_15_15_q ))

	.dataa(!Xd_0__inst_mult_15_14_q ),
	.datab(!Xd_0__inst_mult_15_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_221 ),
	.sharein(Xd_0__inst_mult_15_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_224 ),
	.cout(Xd_0__inst_mult_15_225 ),
	.shareout(Xd_0__inst_mult_15_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_73 (
// Equation(s):
// Xd_0__inst_mult_10_204  = SUM(( !Xd_0__inst_mult_10_14_q  $ (!Xd_0__inst_mult_10_15_q ) ) + ( Xd_0__inst_mult_10_202  ) + ( Xd_0__inst_mult_10_201  ))
// Xd_0__inst_mult_10_205  = CARRY(( !Xd_0__inst_mult_10_14_q  $ (!Xd_0__inst_mult_10_15_q ) ) + ( Xd_0__inst_mult_10_202  ) + ( Xd_0__inst_mult_10_201  ))
// Xd_0__inst_mult_10_206  = SHARE((Xd_0__inst_mult_10_14_q  & Xd_0__inst_mult_10_15_q ))

	.dataa(!Xd_0__inst_mult_10_14_q ),
	.datab(!Xd_0__inst_mult_10_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_201 ),
	.sharein(Xd_0__inst_mult_10_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_204 ),
	.cout(Xd_0__inst_mult_10_205 ),
	.shareout(Xd_0__inst_mult_10_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_77 (
// Equation(s):
// Xd_0__inst_mult_11_208  = SUM(( !Xd_0__inst_mult_11_14_q  $ (!Xd_0__inst_mult_11_15_q ) ) + ( Xd_0__inst_mult_11_206  ) + ( Xd_0__inst_mult_11_205  ))
// Xd_0__inst_mult_11_209  = CARRY(( !Xd_0__inst_mult_11_14_q  $ (!Xd_0__inst_mult_11_15_q ) ) + ( Xd_0__inst_mult_11_206  ) + ( Xd_0__inst_mult_11_205  ))
// Xd_0__inst_mult_11_210  = SHARE((Xd_0__inst_mult_11_14_q  & Xd_0__inst_mult_11_15_q ))

	.dataa(!Xd_0__inst_mult_11_14_q ),
	.datab(!Xd_0__inst_mult_11_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_205 ),
	.sharein(Xd_0__inst_mult_11_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_208 ),
	.cout(Xd_0__inst_mult_11_209 ),
	.shareout(Xd_0__inst_mult_11_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_77 (
// Equation(s):
// Xd_0__inst_mult_8_208  = SUM(( !Xd_0__inst_mult_8_14_q  $ (!Xd_0__inst_mult_8_15_q ) ) + ( Xd_0__inst_mult_8_206  ) + ( Xd_0__inst_mult_8_205  ))
// Xd_0__inst_mult_8_209  = CARRY(( !Xd_0__inst_mult_8_14_q  $ (!Xd_0__inst_mult_8_15_q ) ) + ( Xd_0__inst_mult_8_206  ) + ( Xd_0__inst_mult_8_205  ))
// Xd_0__inst_mult_8_210  = SHARE((Xd_0__inst_mult_8_14_q  & Xd_0__inst_mult_8_15_q ))

	.dataa(!Xd_0__inst_mult_8_14_q ),
	.datab(!Xd_0__inst_mult_8_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_205 ),
	.sharein(Xd_0__inst_mult_8_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_208 ),
	.cout(Xd_0__inst_mult_8_209 ),
	.shareout(Xd_0__inst_mult_8_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_73 (
// Equation(s):
// Xd_0__inst_mult_9_204  = SUM(( !Xd_0__inst_mult_9_14_q  $ (!Xd_0__inst_mult_9_15_q ) ) + ( Xd_0__inst_mult_9_202  ) + ( Xd_0__inst_mult_9_201  ))
// Xd_0__inst_mult_9_205  = CARRY(( !Xd_0__inst_mult_9_14_q  $ (!Xd_0__inst_mult_9_15_q ) ) + ( Xd_0__inst_mult_9_202  ) + ( Xd_0__inst_mult_9_201  ))
// Xd_0__inst_mult_9_206  = SHARE((Xd_0__inst_mult_9_14_q  & Xd_0__inst_mult_9_15_q ))

	.dataa(!Xd_0__inst_mult_9_14_q ),
	.datab(!Xd_0__inst_mult_9_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_201 ),
	.sharein(Xd_0__inst_mult_9_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_204 ),
	.cout(Xd_0__inst_mult_9_205 ),
	.shareout(Xd_0__inst_mult_9_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_73 (
// Equation(s):
// Xd_0__inst_mult_6_204  = SUM(( !Xd_0__inst_mult_6_14_q  $ (!Xd_0__inst_mult_6_15_q ) ) + ( Xd_0__inst_mult_6_202  ) + ( Xd_0__inst_mult_6_201  ))
// Xd_0__inst_mult_6_205  = CARRY(( !Xd_0__inst_mult_6_14_q  $ (!Xd_0__inst_mult_6_15_q ) ) + ( Xd_0__inst_mult_6_202  ) + ( Xd_0__inst_mult_6_201  ))
// Xd_0__inst_mult_6_206  = SHARE((Xd_0__inst_mult_6_14_q  & Xd_0__inst_mult_6_15_q ))

	.dataa(!Xd_0__inst_mult_6_14_q ),
	.datab(!Xd_0__inst_mult_6_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_201 ),
	.sharein(Xd_0__inst_mult_6_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_204 ),
	.cout(Xd_0__inst_mult_6_205 ),
	.shareout(Xd_0__inst_mult_6_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_71 (
// Equation(s):
// Xd_0__inst_mult_7_196  = SUM(( !Xd_0__inst_mult_7_14_q  $ (!Xd_0__inst_mult_7_15_q ) ) + ( Xd_0__inst_mult_7_194  ) + ( Xd_0__inst_mult_7_193  ))
// Xd_0__inst_mult_7_197  = CARRY(( !Xd_0__inst_mult_7_14_q  $ (!Xd_0__inst_mult_7_15_q ) ) + ( Xd_0__inst_mult_7_194  ) + ( Xd_0__inst_mult_7_193  ))
// Xd_0__inst_mult_7_198  = SHARE((Xd_0__inst_mult_7_14_q  & Xd_0__inst_mult_7_15_q ))

	.dataa(!Xd_0__inst_mult_7_14_q ),
	.datab(!Xd_0__inst_mult_7_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_193 ),
	.sharein(Xd_0__inst_mult_7_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_196 ),
	.cout(Xd_0__inst_mult_7_197 ),
	.shareout(Xd_0__inst_mult_7_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_81 (
// Equation(s):
// Xd_0__inst_mult_4_224  = SUM(( !Xd_0__inst_mult_4_14_q  $ (!Xd_0__inst_mult_4_15_q ) ) + ( Xd_0__inst_mult_4_222  ) + ( Xd_0__inst_mult_4_221  ))
// Xd_0__inst_mult_4_225  = CARRY(( !Xd_0__inst_mult_4_14_q  $ (!Xd_0__inst_mult_4_15_q ) ) + ( Xd_0__inst_mult_4_222  ) + ( Xd_0__inst_mult_4_221  ))
// Xd_0__inst_mult_4_226  = SHARE((Xd_0__inst_mult_4_14_q  & Xd_0__inst_mult_4_15_q ))

	.dataa(!Xd_0__inst_mult_4_14_q ),
	.datab(!Xd_0__inst_mult_4_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_221 ),
	.sharein(Xd_0__inst_mult_4_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_224 ),
	.cout(Xd_0__inst_mult_4_225 ),
	.shareout(Xd_0__inst_mult_4_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_71 (
// Equation(s):
// Xd_0__inst_mult_5_196  = SUM(( !Xd_0__inst_mult_5_14_q  $ (!Xd_0__inst_mult_5_15_q ) ) + ( Xd_0__inst_mult_5_194  ) + ( Xd_0__inst_mult_5_193  ))
// Xd_0__inst_mult_5_197  = CARRY(( !Xd_0__inst_mult_5_14_q  $ (!Xd_0__inst_mult_5_15_q ) ) + ( Xd_0__inst_mult_5_194  ) + ( Xd_0__inst_mult_5_193  ))
// Xd_0__inst_mult_5_198  = SHARE((Xd_0__inst_mult_5_14_q  & Xd_0__inst_mult_5_15_q ))

	.dataa(!Xd_0__inst_mult_5_14_q ),
	.datab(!Xd_0__inst_mult_5_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_193 ),
	.sharein(Xd_0__inst_mult_5_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_196 ),
	.cout(Xd_0__inst_mult_5_197 ),
	.shareout(Xd_0__inst_mult_5_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_75 (
// Equation(s):
// Xd_0__inst_mult_2_200  = SUM(( !Xd_0__inst_mult_2_14_q  $ (!Xd_0__inst_mult_2_15_q ) ) + ( Xd_0__inst_mult_2_198  ) + ( Xd_0__inst_mult_2_197  ))
// Xd_0__inst_mult_2_201  = CARRY(( !Xd_0__inst_mult_2_14_q  $ (!Xd_0__inst_mult_2_15_q ) ) + ( Xd_0__inst_mult_2_198  ) + ( Xd_0__inst_mult_2_197  ))
// Xd_0__inst_mult_2_202  = SHARE((Xd_0__inst_mult_2_14_q  & Xd_0__inst_mult_2_15_q ))

	.dataa(!Xd_0__inst_mult_2_14_q ),
	.datab(!Xd_0__inst_mult_2_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_197 ),
	.sharein(Xd_0__inst_mult_2_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_200 ),
	.cout(Xd_0__inst_mult_2_201 ),
	.shareout(Xd_0__inst_mult_2_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_71 (
// Equation(s):
// Xd_0__inst_mult_3_196  = SUM(( !Xd_0__inst_mult_3_14_q  $ (!Xd_0__inst_mult_3_15_q ) ) + ( Xd_0__inst_mult_3_194  ) + ( Xd_0__inst_mult_3_193  ))
// Xd_0__inst_mult_3_197  = CARRY(( !Xd_0__inst_mult_3_14_q  $ (!Xd_0__inst_mult_3_15_q ) ) + ( Xd_0__inst_mult_3_194  ) + ( Xd_0__inst_mult_3_193  ))
// Xd_0__inst_mult_3_198  = SHARE((Xd_0__inst_mult_3_14_q  & Xd_0__inst_mult_3_15_q ))

	.dataa(!Xd_0__inst_mult_3_14_q ),
	.datab(!Xd_0__inst_mult_3_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_193 ),
	.sharein(Xd_0__inst_mult_3_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_196 ),
	.cout(Xd_0__inst_mult_3_197 ),
	.shareout(Xd_0__inst_mult_3_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_75 (
// Equation(s):
// Xd_0__inst_mult_0_200  = SUM(( !Xd_0__inst_mult_0_14_q  $ (!Xd_0__inst_mult_0_15_q ) ) + ( Xd_0__inst_mult_0_198  ) + ( Xd_0__inst_mult_0_197  ))
// Xd_0__inst_mult_0_201  = CARRY(( !Xd_0__inst_mult_0_14_q  $ (!Xd_0__inst_mult_0_15_q ) ) + ( Xd_0__inst_mult_0_198  ) + ( Xd_0__inst_mult_0_197  ))
// Xd_0__inst_mult_0_202  = SHARE((Xd_0__inst_mult_0_14_q  & Xd_0__inst_mult_0_15_q ))

	.dataa(!Xd_0__inst_mult_0_14_q ),
	.datab(!Xd_0__inst_mult_0_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_197 ),
	.sharein(Xd_0__inst_mult_0_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_200 ),
	.cout(Xd_0__inst_mult_0_201 ),
	.shareout(Xd_0__inst_mult_0_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_75 (
// Equation(s):
// Xd_0__inst_mult_1_200  = SUM(( !Xd_0__inst_mult_1_14_q  $ (!Xd_0__inst_mult_1_15_q ) ) + ( Xd_0__inst_mult_1_198  ) + ( Xd_0__inst_mult_1_197  ))
// Xd_0__inst_mult_1_201  = CARRY(( !Xd_0__inst_mult_1_14_q  $ (!Xd_0__inst_mult_1_15_q ) ) + ( Xd_0__inst_mult_1_198  ) + ( Xd_0__inst_mult_1_197  ))
// Xd_0__inst_mult_1_202  = SHARE((Xd_0__inst_mult_1_14_q  & Xd_0__inst_mult_1_15_q ))

	.dataa(!Xd_0__inst_mult_1_14_q ),
	.datab(!Xd_0__inst_mult_1_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_197 ),
	.sharein(Xd_0__inst_mult_1_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_200 ),
	.cout(Xd_0__inst_mult_1_201 ),
	.shareout(Xd_0__inst_mult_1_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_78 (
// Equation(s):
// Xd_0__inst_mult_12_224  = SUM(( !Xd_0__inst_mult_12_16_q  $ (!Xd_0__inst_mult_12_17_q ) ) + ( Xd_0__inst_mult_12_222  ) + ( Xd_0__inst_mult_12_221  ))
// Xd_0__inst_mult_12_225  = CARRY(( !Xd_0__inst_mult_12_16_q  $ (!Xd_0__inst_mult_12_17_q ) ) + ( Xd_0__inst_mult_12_222  ) + ( Xd_0__inst_mult_12_221  ))
// Xd_0__inst_mult_12_226  = SHARE((Xd_0__inst_mult_12_16_q  & Xd_0__inst_mult_12_17_q ))

	.dataa(!Xd_0__inst_mult_12_16_q ),
	.datab(!Xd_0__inst_mult_12_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_221 ),
	.sharein(Xd_0__inst_mult_12_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_224 ),
	.cout(Xd_0__inst_mult_12_225 ),
	.shareout(Xd_0__inst_mult_12_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_78 (
// Equation(s):
// Xd_0__inst_mult_13_212  = SUM(( !Xd_0__inst_mult_13_16_q  $ (!Xd_0__inst_mult_13_17_q ) ) + ( Xd_0__inst_mult_13_210  ) + ( Xd_0__inst_mult_13_209  ))
// Xd_0__inst_mult_13_213  = CARRY(( !Xd_0__inst_mult_13_16_q  $ (!Xd_0__inst_mult_13_17_q ) ) + ( Xd_0__inst_mult_13_210  ) + ( Xd_0__inst_mult_13_209  ))
// Xd_0__inst_mult_13_214  = SHARE((Xd_0__inst_mult_13_16_q  & Xd_0__inst_mult_13_17_q ))

	.dataa(!Xd_0__inst_mult_13_16_q ),
	.datab(!Xd_0__inst_mult_13_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_209 ),
	.sharein(Xd_0__inst_mult_13_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_212 ),
	.cout(Xd_0__inst_mult_13_213 ),
	.shareout(Xd_0__inst_mult_13_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_82 (
// Equation(s):
// Xd_0__inst_mult_14_228  = SUM(( !Xd_0__inst_mult_14_16_q  $ (!Xd_0__inst_mult_14_17_q ) ) + ( Xd_0__inst_mult_14_226  ) + ( Xd_0__inst_mult_14_225  ))
// Xd_0__inst_mult_14_229  = CARRY(( !Xd_0__inst_mult_14_16_q  $ (!Xd_0__inst_mult_14_17_q ) ) + ( Xd_0__inst_mult_14_226  ) + ( Xd_0__inst_mult_14_225  ))
// Xd_0__inst_mult_14_230  = SHARE((Xd_0__inst_mult_14_16_q  & Xd_0__inst_mult_14_17_q ))

	.dataa(!Xd_0__inst_mult_14_16_q ),
	.datab(!Xd_0__inst_mult_14_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_225 ),
	.sharein(Xd_0__inst_mult_14_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_228 ),
	.cout(Xd_0__inst_mult_14_229 ),
	.shareout(Xd_0__inst_mult_14_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_82 (
// Equation(s):
// Xd_0__inst_mult_15_228  = SUM(( !Xd_0__inst_mult_15_16_q  $ (!Xd_0__inst_mult_15_17_q ) ) + ( Xd_0__inst_mult_15_226  ) + ( Xd_0__inst_mult_15_225  ))
// Xd_0__inst_mult_15_229  = CARRY(( !Xd_0__inst_mult_15_16_q  $ (!Xd_0__inst_mult_15_17_q ) ) + ( Xd_0__inst_mult_15_226  ) + ( Xd_0__inst_mult_15_225  ))
// Xd_0__inst_mult_15_230  = SHARE((Xd_0__inst_mult_15_16_q  & Xd_0__inst_mult_15_17_q ))

	.dataa(!Xd_0__inst_mult_15_16_q ),
	.datab(!Xd_0__inst_mult_15_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_225 ),
	.sharein(Xd_0__inst_mult_15_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_228 ),
	.cout(Xd_0__inst_mult_15_229 ),
	.shareout(Xd_0__inst_mult_15_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_74 (
// Equation(s):
// Xd_0__inst_mult_10_208  = SUM(( !Xd_0__inst_mult_10_16_q  $ (!Xd_0__inst_mult_10_17_q ) ) + ( Xd_0__inst_mult_10_206  ) + ( Xd_0__inst_mult_10_205  ))
// Xd_0__inst_mult_10_209  = CARRY(( !Xd_0__inst_mult_10_16_q  $ (!Xd_0__inst_mult_10_17_q ) ) + ( Xd_0__inst_mult_10_206  ) + ( Xd_0__inst_mult_10_205  ))
// Xd_0__inst_mult_10_210  = SHARE((Xd_0__inst_mult_10_16_q  & Xd_0__inst_mult_10_17_q ))

	.dataa(!Xd_0__inst_mult_10_16_q ),
	.datab(!Xd_0__inst_mult_10_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_205 ),
	.sharein(Xd_0__inst_mult_10_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_208 ),
	.cout(Xd_0__inst_mult_10_209 ),
	.shareout(Xd_0__inst_mult_10_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_78 (
// Equation(s):
// Xd_0__inst_mult_11_212  = SUM(( !Xd_0__inst_mult_11_16_q  $ (!Xd_0__inst_mult_11_17_q ) ) + ( Xd_0__inst_mult_11_210  ) + ( Xd_0__inst_mult_11_209  ))
// Xd_0__inst_mult_11_213  = CARRY(( !Xd_0__inst_mult_11_16_q  $ (!Xd_0__inst_mult_11_17_q ) ) + ( Xd_0__inst_mult_11_210  ) + ( Xd_0__inst_mult_11_209  ))
// Xd_0__inst_mult_11_214  = SHARE((Xd_0__inst_mult_11_16_q  & Xd_0__inst_mult_11_17_q ))

	.dataa(!Xd_0__inst_mult_11_16_q ),
	.datab(!Xd_0__inst_mult_11_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_209 ),
	.sharein(Xd_0__inst_mult_11_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_212 ),
	.cout(Xd_0__inst_mult_11_213 ),
	.shareout(Xd_0__inst_mult_11_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_78 (
// Equation(s):
// Xd_0__inst_mult_8_212  = SUM(( !Xd_0__inst_mult_8_16_q  $ (!Xd_0__inst_mult_8_17_q ) ) + ( Xd_0__inst_mult_8_210  ) + ( Xd_0__inst_mult_8_209  ))
// Xd_0__inst_mult_8_213  = CARRY(( !Xd_0__inst_mult_8_16_q  $ (!Xd_0__inst_mult_8_17_q ) ) + ( Xd_0__inst_mult_8_210  ) + ( Xd_0__inst_mult_8_209  ))
// Xd_0__inst_mult_8_214  = SHARE((Xd_0__inst_mult_8_16_q  & Xd_0__inst_mult_8_17_q ))

	.dataa(!Xd_0__inst_mult_8_16_q ),
	.datab(!Xd_0__inst_mult_8_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_209 ),
	.sharein(Xd_0__inst_mult_8_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_212 ),
	.cout(Xd_0__inst_mult_8_213 ),
	.shareout(Xd_0__inst_mult_8_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_74 (
// Equation(s):
// Xd_0__inst_mult_9_208  = SUM(( !Xd_0__inst_mult_9_16_q  $ (!Xd_0__inst_mult_9_17_q ) ) + ( Xd_0__inst_mult_9_206  ) + ( Xd_0__inst_mult_9_205  ))
// Xd_0__inst_mult_9_209  = CARRY(( !Xd_0__inst_mult_9_16_q  $ (!Xd_0__inst_mult_9_17_q ) ) + ( Xd_0__inst_mult_9_206  ) + ( Xd_0__inst_mult_9_205  ))
// Xd_0__inst_mult_9_210  = SHARE((Xd_0__inst_mult_9_16_q  & Xd_0__inst_mult_9_17_q ))

	.dataa(!Xd_0__inst_mult_9_16_q ),
	.datab(!Xd_0__inst_mult_9_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_205 ),
	.sharein(Xd_0__inst_mult_9_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_208 ),
	.cout(Xd_0__inst_mult_9_209 ),
	.shareout(Xd_0__inst_mult_9_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_74 (
// Equation(s):
// Xd_0__inst_mult_6_208  = SUM(( !Xd_0__inst_mult_6_16_q  $ (!Xd_0__inst_mult_6_17_q ) ) + ( Xd_0__inst_mult_6_206  ) + ( Xd_0__inst_mult_6_205  ))
// Xd_0__inst_mult_6_209  = CARRY(( !Xd_0__inst_mult_6_16_q  $ (!Xd_0__inst_mult_6_17_q ) ) + ( Xd_0__inst_mult_6_206  ) + ( Xd_0__inst_mult_6_205  ))
// Xd_0__inst_mult_6_210  = SHARE((Xd_0__inst_mult_6_16_q  & Xd_0__inst_mult_6_17_q ))

	.dataa(!Xd_0__inst_mult_6_16_q ),
	.datab(!Xd_0__inst_mult_6_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_205 ),
	.sharein(Xd_0__inst_mult_6_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_208 ),
	.cout(Xd_0__inst_mult_6_209 ),
	.shareout(Xd_0__inst_mult_6_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_72 (
// Equation(s):
// Xd_0__inst_mult_7_200  = SUM(( !Xd_0__inst_mult_7_16_q  $ (!Xd_0__inst_mult_7_17_q ) ) + ( Xd_0__inst_mult_7_198  ) + ( Xd_0__inst_mult_7_197  ))
// Xd_0__inst_mult_7_201  = CARRY(( !Xd_0__inst_mult_7_16_q  $ (!Xd_0__inst_mult_7_17_q ) ) + ( Xd_0__inst_mult_7_198  ) + ( Xd_0__inst_mult_7_197  ))
// Xd_0__inst_mult_7_202  = SHARE((Xd_0__inst_mult_7_16_q  & Xd_0__inst_mult_7_17_q ))

	.dataa(!Xd_0__inst_mult_7_16_q ),
	.datab(!Xd_0__inst_mult_7_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_197 ),
	.sharein(Xd_0__inst_mult_7_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_200 ),
	.cout(Xd_0__inst_mult_7_201 ),
	.shareout(Xd_0__inst_mult_7_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_82 (
// Equation(s):
// Xd_0__inst_mult_4_228  = SUM(( !Xd_0__inst_mult_4_16_q  $ (!Xd_0__inst_mult_4_17_q ) ) + ( Xd_0__inst_mult_4_226  ) + ( Xd_0__inst_mult_4_225  ))
// Xd_0__inst_mult_4_229  = CARRY(( !Xd_0__inst_mult_4_16_q  $ (!Xd_0__inst_mult_4_17_q ) ) + ( Xd_0__inst_mult_4_226  ) + ( Xd_0__inst_mult_4_225  ))
// Xd_0__inst_mult_4_230  = SHARE((Xd_0__inst_mult_4_16_q  & Xd_0__inst_mult_4_17_q ))

	.dataa(!Xd_0__inst_mult_4_16_q ),
	.datab(!Xd_0__inst_mult_4_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_225 ),
	.sharein(Xd_0__inst_mult_4_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_228 ),
	.cout(Xd_0__inst_mult_4_229 ),
	.shareout(Xd_0__inst_mult_4_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_72 (
// Equation(s):
// Xd_0__inst_mult_5_200  = SUM(( !Xd_0__inst_mult_5_16_q  $ (!Xd_0__inst_mult_5_17_q ) ) + ( Xd_0__inst_mult_5_198  ) + ( Xd_0__inst_mult_5_197  ))
// Xd_0__inst_mult_5_201  = CARRY(( !Xd_0__inst_mult_5_16_q  $ (!Xd_0__inst_mult_5_17_q ) ) + ( Xd_0__inst_mult_5_198  ) + ( Xd_0__inst_mult_5_197  ))
// Xd_0__inst_mult_5_202  = SHARE((Xd_0__inst_mult_5_16_q  & Xd_0__inst_mult_5_17_q ))

	.dataa(!Xd_0__inst_mult_5_16_q ),
	.datab(!Xd_0__inst_mult_5_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_197 ),
	.sharein(Xd_0__inst_mult_5_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_200 ),
	.cout(Xd_0__inst_mult_5_201 ),
	.shareout(Xd_0__inst_mult_5_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_76 (
// Equation(s):
// Xd_0__inst_mult_2_204  = SUM(( !Xd_0__inst_mult_2_16_q  $ (!Xd_0__inst_mult_2_17_q ) ) + ( Xd_0__inst_mult_2_202  ) + ( Xd_0__inst_mult_2_201  ))
// Xd_0__inst_mult_2_205  = CARRY(( !Xd_0__inst_mult_2_16_q  $ (!Xd_0__inst_mult_2_17_q ) ) + ( Xd_0__inst_mult_2_202  ) + ( Xd_0__inst_mult_2_201  ))
// Xd_0__inst_mult_2_206  = SHARE((Xd_0__inst_mult_2_16_q  & Xd_0__inst_mult_2_17_q ))

	.dataa(!Xd_0__inst_mult_2_16_q ),
	.datab(!Xd_0__inst_mult_2_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_201 ),
	.sharein(Xd_0__inst_mult_2_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_204 ),
	.cout(Xd_0__inst_mult_2_205 ),
	.shareout(Xd_0__inst_mult_2_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_72 (
// Equation(s):
// Xd_0__inst_mult_3_200  = SUM(( !Xd_0__inst_mult_3_16_q  $ (!Xd_0__inst_mult_3_17_q ) ) + ( Xd_0__inst_mult_3_198  ) + ( Xd_0__inst_mult_3_197  ))
// Xd_0__inst_mult_3_201  = CARRY(( !Xd_0__inst_mult_3_16_q  $ (!Xd_0__inst_mult_3_17_q ) ) + ( Xd_0__inst_mult_3_198  ) + ( Xd_0__inst_mult_3_197  ))
// Xd_0__inst_mult_3_202  = SHARE((Xd_0__inst_mult_3_16_q  & Xd_0__inst_mult_3_17_q ))

	.dataa(!Xd_0__inst_mult_3_16_q ),
	.datab(!Xd_0__inst_mult_3_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_197 ),
	.sharein(Xd_0__inst_mult_3_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_200 ),
	.cout(Xd_0__inst_mult_3_201 ),
	.shareout(Xd_0__inst_mult_3_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_76 (
// Equation(s):
// Xd_0__inst_mult_0_204  = SUM(( !Xd_0__inst_mult_0_16_q  $ (!Xd_0__inst_mult_0_17_q ) ) + ( Xd_0__inst_mult_0_202  ) + ( Xd_0__inst_mult_0_201  ))
// Xd_0__inst_mult_0_205  = CARRY(( !Xd_0__inst_mult_0_16_q  $ (!Xd_0__inst_mult_0_17_q ) ) + ( Xd_0__inst_mult_0_202  ) + ( Xd_0__inst_mult_0_201  ))
// Xd_0__inst_mult_0_206  = SHARE((Xd_0__inst_mult_0_16_q  & Xd_0__inst_mult_0_17_q ))

	.dataa(!Xd_0__inst_mult_0_16_q ),
	.datab(!Xd_0__inst_mult_0_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_201 ),
	.sharein(Xd_0__inst_mult_0_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_204 ),
	.cout(Xd_0__inst_mult_0_205 ),
	.shareout(Xd_0__inst_mult_0_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_76 (
// Equation(s):
// Xd_0__inst_mult_1_204  = SUM(( !Xd_0__inst_mult_1_16_q  $ (!Xd_0__inst_mult_1_17_q ) ) + ( Xd_0__inst_mult_1_202  ) + ( Xd_0__inst_mult_1_201  ))
// Xd_0__inst_mult_1_205  = CARRY(( !Xd_0__inst_mult_1_16_q  $ (!Xd_0__inst_mult_1_17_q ) ) + ( Xd_0__inst_mult_1_202  ) + ( Xd_0__inst_mult_1_201  ))
// Xd_0__inst_mult_1_206  = SHARE((Xd_0__inst_mult_1_16_q  & Xd_0__inst_mult_1_17_q ))

	.dataa(!Xd_0__inst_mult_1_16_q ),
	.datab(!Xd_0__inst_mult_1_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_201 ),
	.sharein(Xd_0__inst_mult_1_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_204 ),
	.cout(Xd_0__inst_mult_1_205 ),
	.shareout(Xd_0__inst_mult_1_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_79 (
// Equation(s):
// Xd_0__inst_mult_12_228  = SUM(( !Xd_0__inst_mult_12_18_q  $ (!Xd_0__inst_mult_12_19_q ) ) + ( Xd_0__inst_mult_12_226  ) + ( Xd_0__inst_mult_12_225  ))
// Xd_0__inst_mult_12_229  = CARRY(( !Xd_0__inst_mult_12_18_q  $ (!Xd_0__inst_mult_12_19_q ) ) + ( Xd_0__inst_mult_12_226  ) + ( Xd_0__inst_mult_12_225  ))
// Xd_0__inst_mult_12_230  = SHARE((Xd_0__inst_mult_12_18_q  & Xd_0__inst_mult_12_19_q ))

	.dataa(!Xd_0__inst_mult_12_18_q ),
	.datab(!Xd_0__inst_mult_12_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_225 ),
	.sharein(Xd_0__inst_mult_12_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_228 ),
	.cout(Xd_0__inst_mult_12_229 ),
	.shareout(Xd_0__inst_mult_12_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_79 (
// Equation(s):
// Xd_0__inst_mult_13_216  = SUM(( !Xd_0__inst_mult_13_18_q  $ (!Xd_0__inst_mult_13_19_q ) ) + ( Xd_0__inst_mult_13_214  ) + ( Xd_0__inst_mult_13_213  ))
// Xd_0__inst_mult_13_217  = CARRY(( !Xd_0__inst_mult_13_18_q  $ (!Xd_0__inst_mult_13_19_q ) ) + ( Xd_0__inst_mult_13_214  ) + ( Xd_0__inst_mult_13_213  ))
// Xd_0__inst_mult_13_218  = SHARE((Xd_0__inst_mult_13_18_q  & Xd_0__inst_mult_13_19_q ))

	.dataa(!Xd_0__inst_mult_13_18_q ),
	.datab(!Xd_0__inst_mult_13_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_213 ),
	.sharein(Xd_0__inst_mult_13_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_216 ),
	.cout(Xd_0__inst_mult_13_217 ),
	.shareout(Xd_0__inst_mult_13_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_83 (
// Equation(s):
// Xd_0__inst_mult_14_232  = SUM(( !Xd_0__inst_mult_14_18_q  $ (!Xd_0__inst_mult_14_19_q ) ) + ( Xd_0__inst_mult_14_230  ) + ( Xd_0__inst_mult_14_229  ))
// Xd_0__inst_mult_14_233  = CARRY(( !Xd_0__inst_mult_14_18_q  $ (!Xd_0__inst_mult_14_19_q ) ) + ( Xd_0__inst_mult_14_230  ) + ( Xd_0__inst_mult_14_229  ))
// Xd_0__inst_mult_14_234  = SHARE((Xd_0__inst_mult_14_18_q  & Xd_0__inst_mult_14_19_q ))

	.dataa(!Xd_0__inst_mult_14_18_q ),
	.datab(!Xd_0__inst_mult_14_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_229 ),
	.sharein(Xd_0__inst_mult_14_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_232 ),
	.cout(Xd_0__inst_mult_14_233 ),
	.shareout(Xd_0__inst_mult_14_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_83 (
// Equation(s):
// Xd_0__inst_mult_15_232  = SUM(( !Xd_0__inst_mult_15_18_q  $ (!Xd_0__inst_mult_15_19_q ) ) + ( Xd_0__inst_mult_15_230  ) + ( Xd_0__inst_mult_15_229  ))
// Xd_0__inst_mult_15_233  = CARRY(( !Xd_0__inst_mult_15_18_q  $ (!Xd_0__inst_mult_15_19_q ) ) + ( Xd_0__inst_mult_15_230  ) + ( Xd_0__inst_mult_15_229  ))
// Xd_0__inst_mult_15_234  = SHARE((Xd_0__inst_mult_15_18_q  & Xd_0__inst_mult_15_19_q ))

	.dataa(!Xd_0__inst_mult_15_18_q ),
	.datab(!Xd_0__inst_mult_15_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_229 ),
	.sharein(Xd_0__inst_mult_15_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_232 ),
	.cout(Xd_0__inst_mult_15_233 ),
	.shareout(Xd_0__inst_mult_15_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_75 (
// Equation(s):
// Xd_0__inst_mult_10_212  = SUM(( !Xd_0__inst_mult_10_18_q  $ (!Xd_0__inst_mult_10_19_q ) ) + ( Xd_0__inst_mult_10_210  ) + ( Xd_0__inst_mult_10_209  ))
// Xd_0__inst_mult_10_213  = CARRY(( !Xd_0__inst_mult_10_18_q  $ (!Xd_0__inst_mult_10_19_q ) ) + ( Xd_0__inst_mult_10_210  ) + ( Xd_0__inst_mult_10_209  ))
// Xd_0__inst_mult_10_214  = SHARE((Xd_0__inst_mult_10_18_q  & Xd_0__inst_mult_10_19_q ))

	.dataa(!Xd_0__inst_mult_10_18_q ),
	.datab(!Xd_0__inst_mult_10_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_209 ),
	.sharein(Xd_0__inst_mult_10_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_212 ),
	.cout(Xd_0__inst_mult_10_213 ),
	.shareout(Xd_0__inst_mult_10_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_79 (
// Equation(s):
// Xd_0__inst_mult_11_216  = SUM(( !Xd_0__inst_mult_11_18_q  $ (!Xd_0__inst_mult_11_19_q ) ) + ( Xd_0__inst_mult_11_214  ) + ( Xd_0__inst_mult_11_213  ))
// Xd_0__inst_mult_11_217  = CARRY(( !Xd_0__inst_mult_11_18_q  $ (!Xd_0__inst_mult_11_19_q ) ) + ( Xd_0__inst_mult_11_214  ) + ( Xd_0__inst_mult_11_213  ))
// Xd_0__inst_mult_11_218  = SHARE((Xd_0__inst_mult_11_18_q  & Xd_0__inst_mult_11_19_q ))

	.dataa(!Xd_0__inst_mult_11_18_q ),
	.datab(!Xd_0__inst_mult_11_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_213 ),
	.sharein(Xd_0__inst_mult_11_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_216 ),
	.cout(Xd_0__inst_mult_11_217 ),
	.shareout(Xd_0__inst_mult_11_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_79 (
// Equation(s):
// Xd_0__inst_mult_8_216  = SUM(( !Xd_0__inst_mult_8_18_q  $ (!Xd_0__inst_mult_8_19_q ) ) + ( Xd_0__inst_mult_8_214  ) + ( Xd_0__inst_mult_8_213  ))
// Xd_0__inst_mult_8_217  = CARRY(( !Xd_0__inst_mult_8_18_q  $ (!Xd_0__inst_mult_8_19_q ) ) + ( Xd_0__inst_mult_8_214  ) + ( Xd_0__inst_mult_8_213  ))
// Xd_0__inst_mult_8_218  = SHARE((Xd_0__inst_mult_8_18_q  & Xd_0__inst_mult_8_19_q ))

	.dataa(!Xd_0__inst_mult_8_18_q ),
	.datab(!Xd_0__inst_mult_8_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_213 ),
	.sharein(Xd_0__inst_mult_8_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_216 ),
	.cout(Xd_0__inst_mult_8_217 ),
	.shareout(Xd_0__inst_mult_8_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_75 (
// Equation(s):
// Xd_0__inst_mult_9_212  = SUM(( !Xd_0__inst_mult_9_18_q  $ (!Xd_0__inst_mult_9_19_q ) ) + ( Xd_0__inst_mult_9_210  ) + ( Xd_0__inst_mult_9_209  ))
// Xd_0__inst_mult_9_213  = CARRY(( !Xd_0__inst_mult_9_18_q  $ (!Xd_0__inst_mult_9_19_q ) ) + ( Xd_0__inst_mult_9_210  ) + ( Xd_0__inst_mult_9_209  ))
// Xd_0__inst_mult_9_214  = SHARE((Xd_0__inst_mult_9_18_q  & Xd_0__inst_mult_9_19_q ))

	.dataa(!Xd_0__inst_mult_9_18_q ),
	.datab(!Xd_0__inst_mult_9_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_209 ),
	.sharein(Xd_0__inst_mult_9_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_212 ),
	.cout(Xd_0__inst_mult_9_213 ),
	.shareout(Xd_0__inst_mult_9_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_75 (
// Equation(s):
// Xd_0__inst_mult_6_212  = SUM(( !Xd_0__inst_mult_6_18_q  $ (!Xd_0__inst_mult_6_19_q ) ) + ( Xd_0__inst_mult_6_210  ) + ( Xd_0__inst_mult_6_209  ))
// Xd_0__inst_mult_6_213  = CARRY(( !Xd_0__inst_mult_6_18_q  $ (!Xd_0__inst_mult_6_19_q ) ) + ( Xd_0__inst_mult_6_210  ) + ( Xd_0__inst_mult_6_209  ))
// Xd_0__inst_mult_6_214  = SHARE((Xd_0__inst_mult_6_18_q  & Xd_0__inst_mult_6_19_q ))

	.dataa(!Xd_0__inst_mult_6_18_q ),
	.datab(!Xd_0__inst_mult_6_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_209 ),
	.sharein(Xd_0__inst_mult_6_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_212 ),
	.cout(Xd_0__inst_mult_6_213 ),
	.shareout(Xd_0__inst_mult_6_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_73 (
// Equation(s):
// Xd_0__inst_mult_7_204  = SUM(( !Xd_0__inst_mult_7_18_q  $ (!Xd_0__inst_mult_7_19_q ) ) + ( Xd_0__inst_mult_7_202  ) + ( Xd_0__inst_mult_7_201  ))
// Xd_0__inst_mult_7_205  = CARRY(( !Xd_0__inst_mult_7_18_q  $ (!Xd_0__inst_mult_7_19_q ) ) + ( Xd_0__inst_mult_7_202  ) + ( Xd_0__inst_mult_7_201  ))
// Xd_0__inst_mult_7_206  = SHARE((Xd_0__inst_mult_7_18_q  & Xd_0__inst_mult_7_19_q ))

	.dataa(!Xd_0__inst_mult_7_18_q ),
	.datab(!Xd_0__inst_mult_7_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_201 ),
	.sharein(Xd_0__inst_mult_7_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_204 ),
	.cout(Xd_0__inst_mult_7_205 ),
	.shareout(Xd_0__inst_mult_7_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_83 (
// Equation(s):
// Xd_0__inst_mult_4_232  = SUM(( !Xd_0__inst_mult_4_18_q  $ (!Xd_0__inst_mult_4_19_q ) ) + ( Xd_0__inst_mult_4_230  ) + ( Xd_0__inst_mult_4_229  ))
// Xd_0__inst_mult_4_233  = CARRY(( !Xd_0__inst_mult_4_18_q  $ (!Xd_0__inst_mult_4_19_q ) ) + ( Xd_0__inst_mult_4_230  ) + ( Xd_0__inst_mult_4_229  ))
// Xd_0__inst_mult_4_234  = SHARE((Xd_0__inst_mult_4_18_q  & Xd_0__inst_mult_4_19_q ))

	.dataa(!Xd_0__inst_mult_4_18_q ),
	.datab(!Xd_0__inst_mult_4_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_229 ),
	.sharein(Xd_0__inst_mult_4_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_232 ),
	.cout(Xd_0__inst_mult_4_233 ),
	.shareout(Xd_0__inst_mult_4_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_73 (
// Equation(s):
// Xd_0__inst_mult_5_204  = SUM(( !Xd_0__inst_mult_5_18_q  $ (!Xd_0__inst_mult_5_19_q ) ) + ( Xd_0__inst_mult_5_202  ) + ( Xd_0__inst_mult_5_201  ))
// Xd_0__inst_mult_5_205  = CARRY(( !Xd_0__inst_mult_5_18_q  $ (!Xd_0__inst_mult_5_19_q ) ) + ( Xd_0__inst_mult_5_202  ) + ( Xd_0__inst_mult_5_201  ))
// Xd_0__inst_mult_5_206  = SHARE((Xd_0__inst_mult_5_18_q  & Xd_0__inst_mult_5_19_q ))

	.dataa(!Xd_0__inst_mult_5_18_q ),
	.datab(!Xd_0__inst_mult_5_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_201 ),
	.sharein(Xd_0__inst_mult_5_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_204 ),
	.cout(Xd_0__inst_mult_5_205 ),
	.shareout(Xd_0__inst_mult_5_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_77 (
// Equation(s):
// Xd_0__inst_mult_2_208  = SUM(( !Xd_0__inst_mult_2_18_q  $ (!Xd_0__inst_mult_2_19_q ) ) + ( Xd_0__inst_mult_2_206  ) + ( Xd_0__inst_mult_2_205  ))
// Xd_0__inst_mult_2_209  = CARRY(( !Xd_0__inst_mult_2_18_q  $ (!Xd_0__inst_mult_2_19_q ) ) + ( Xd_0__inst_mult_2_206  ) + ( Xd_0__inst_mult_2_205  ))
// Xd_0__inst_mult_2_210  = SHARE((Xd_0__inst_mult_2_18_q  & Xd_0__inst_mult_2_19_q ))

	.dataa(!Xd_0__inst_mult_2_18_q ),
	.datab(!Xd_0__inst_mult_2_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_205 ),
	.sharein(Xd_0__inst_mult_2_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_208 ),
	.cout(Xd_0__inst_mult_2_209 ),
	.shareout(Xd_0__inst_mult_2_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_73 (
// Equation(s):
// Xd_0__inst_mult_3_204  = SUM(( !Xd_0__inst_mult_3_18_q  $ (!Xd_0__inst_mult_3_19_q ) ) + ( Xd_0__inst_mult_3_202  ) + ( Xd_0__inst_mult_3_201  ))
// Xd_0__inst_mult_3_205  = CARRY(( !Xd_0__inst_mult_3_18_q  $ (!Xd_0__inst_mult_3_19_q ) ) + ( Xd_0__inst_mult_3_202  ) + ( Xd_0__inst_mult_3_201  ))
// Xd_0__inst_mult_3_206  = SHARE((Xd_0__inst_mult_3_18_q  & Xd_0__inst_mult_3_19_q ))

	.dataa(!Xd_0__inst_mult_3_18_q ),
	.datab(!Xd_0__inst_mult_3_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_201 ),
	.sharein(Xd_0__inst_mult_3_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_204 ),
	.cout(Xd_0__inst_mult_3_205 ),
	.shareout(Xd_0__inst_mult_3_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_77 (
// Equation(s):
// Xd_0__inst_mult_0_208  = SUM(( !Xd_0__inst_mult_0_18_q  $ (!Xd_0__inst_mult_0_19_q ) ) + ( Xd_0__inst_mult_0_206  ) + ( Xd_0__inst_mult_0_205  ))
// Xd_0__inst_mult_0_209  = CARRY(( !Xd_0__inst_mult_0_18_q  $ (!Xd_0__inst_mult_0_19_q ) ) + ( Xd_0__inst_mult_0_206  ) + ( Xd_0__inst_mult_0_205  ))
// Xd_0__inst_mult_0_210  = SHARE((Xd_0__inst_mult_0_18_q  & Xd_0__inst_mult_0_19_q ))

	.dataa(!Xd_0__inst_mult_0_18_q ),
	.datab(!Xd_0__inst_mult_0_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_205 ),
	.sharein(Xd_0__inst_mult_0_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_208 ),
	.cout(Xd_0__inst_mult_0_209 ),
	.shareout(Xd_0__inst_mult_0_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_77 (
// Equation(s):
// Xd_0__inst_mult_1_208  = SUM(( !Xd_0__inst_mult_1_18_q  $ (!Xd_0__inst_mult_1_19_q ) ) + ( Xd_0__inst_mult_1_206  ) + ( Xd_0__inst_mult_1_205  ))
// Xd_0__inst_mult_1_209  = CARRY(( !Xd_0__inst_mult_1_18_q  $ (!Xd_0__inst_mult_1_19_q ) ) + ( Xd_0__inst_mult_1_206  ) + ( Xd_0__inst_mult_1_205  ))
// Xd_0__inst_mult_1_210  = SHARE((Xd_0__inst_mult_1_18_q  & Xd_0__inst_mult_1_19_q ))

	.dataa(!Xd_0__inst_mult_1_18_q ),
	.datab(!Xd_0__inst_mult_1_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_205 ),
	.sharein(Xd_0__inst_mult_1_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_208 ),
	.cout(Xd_0__inst_mult_1_209 ),
	.shareout(Xd_0__inst_mult_1_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_80 (
// Equation(s):
// Xd_0__inst_mult_12_232  = SUM(( !Xd_0__inst_mult_12_20_q  $ (!Xd_0__inst_mult_12_21_q  $ (((Xd_0__inst_mult_12_22_q  & Xd_0__inst_mult_12_23_q )))) ) + ( Xd_0__inst_mult_12_230  ) + ( Xd_0__inst_mult_12_229  ))
// Xd_0__inst_mult_12_233  = CARRY(( !Xd_0__inst_mult_12_20_q  $ (!Xd_0__inst_mult_12_21_q  $ (((Xd_0__inst_mult_12_22_q  & Xd_0__inst_mult_12_23_q )))) ) + ( Xd_0__inst_mult_12_230  ) + ( Xd_0__inst_mult_12_229  ))
// Xd_0__inst_mult_12_234  = SHARE((Xd_0__inst_mult_12_22_q  & (Xd_0__inst_mult_12_23_q  & (!Xd_0__inst_mult_12_20_q  $ (!Xd_0__inst_mult_12_21_q )))))

	.dataa(!Xd_0__inst_mult_12_20_q ),
	.datab(!Xd_0__inst_mult_12_21_q ),
	.datac(!Xd_0__inst_mult_12_22_q ),
	.datad(!Xd_0__inst_mult_12_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_229 ),
	.sharein(Xd_0__inst_mult_12_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_232 ),
	.cout(Xd_0__inst_mult_12_233 ),
	.shareout(Xd_0__inst_mult_12_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_80 (
// Equation(s):
// Xd_0__inst_mult_13_220  = SUM(( !Xd_0__inst_mult_13_20_q  $ (!Xd_0__inst_mult_13_21_q  $ (((Xd_0__inst_mult_13_22_q  & Xd_0__inst_mult_13_23_q )))) ) + ( Xd_0__inst_mult_13_218  ) + ( Xd_0__inst_mult_13_217  ))
// Xd_0__inst_mult_13_221  = CARRY(( !Xd_0__inst_mult_13_20_q  $ (!Xd_0__inst_mult_13_21_q  $ (((Xd_0__inst_mult_13_22_q  & Xd_0__inst_mult_13_23_q )))) ) + ( Xd_0__inst_mult_13_218  ) + ( Xd_0__inst_mult_13_217  ))
// Xd_0__inst_mult_13_222  = SHARE((Xd_0__inst_mult_13_22_q  & (Xd_0__inst_mult_13_23_q  & (!Xd_0__inst_mult_13_20_q  $ (!Xd_0__inst_mult_13_21_q )))))

	.dataa(!Xd_0__inst_mult_13_20_q ),
	.datab(!Xd_0__inst_mult_13_21_q ),
	.datac(!Xd_0__inst_mult_13_22_q ),
	.datad(!Xd_0__inst_mult_13_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_217 ),
	.sharein(Xd_0__inst_mult_13_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_220 ),
	.cout(Xd_0__inst_mult_13_221 ),
	.shareout(Xd_0__inst_mult_13_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_84 (
// Equation(s):
// Xd_0__inst_mult_14_236  = SUM(( !Xd_0__inst_mult_14_20_q  $ (!Xd_0__inst_mult_14_21_q  $ (((Xd_0__inst_mult_14_22_q  & Xd_0__inst_mult_14_23_q )))) ) + ( Xd_0__inst_mult_14_234  ) + ( Xd_0__inst_mult_14_233  ))
// Xd_0__inst_mult_14_237  = CARRY(( !Xd_0__inst_mult_14_20_q  $ (!Xd_0__inst_mult_14_21_q  $ (((Xd_0__inst_mult_14_22_q  & Xd_0__inst_mult_14_23_q )))) ) + ( Xd_0__inst_mult_14_234  ) + ( Xd_0__inst_mult_14_233  ))
// Xd_0__inst_mult_14_238  = SHARE((Xd_0__inst_mult_14_22_q  & (Xd_0__inst_mult_14_23_q  & (!Xd_0__inst_mult_14_20_q  $ (!Xd_0__inst_mult_14_21_q )))))

	.dataa(!Xd_0__inst_mult_14_20_q ),
	.datab(!Xd_0__inst_mult_14_21_q ),
	.datac(!Xd_0__inst_mult_14_22_q ),
	.datad(!Xd_0__inst_mult_14_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_233 ),
	.sharein(Xd_0__inst_mult_14_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_236 ),
	.cout(Xd_0__inst_mult_14_237 ),
	.shareout(Xd_0__inst_mult_14_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_84 (
// Equation(s):
// Xd_0__inst_mult_15_236  = SUM(( !Xd_0__inst_mult_15_20_q  $ (!Xd_0__inst_mult_15_21_q  $ (((Xd_0__inst_mult_15_22_q  & Xd_0__inst_mult_15_23_q )))) ) + ( Xd_0__inst_mult_15_234  ) + ( Xd_0__inst_mult_15_233  ))
// Xd_0__inst_mult_15_237  = CARRY(( !Xd_0__inst_mult_15_20_q  $ (!Xd_0__inst_mult_15_21_q  $ (((Xd_0__inst_mult_15_22_q  & Xd_0__inst_mult_15_23_q )))) ) + ( Xd_0__inst_mult_15_234  ) + ( Xd_0__inst_mult_15_233  ))
// Xd_0__inst_mult_15_238  = SHARE((Xd_0__inst_mult_15_22_q  & (Xd_0__inst_mult_15_23_q  & (!Xd_0__inst_mult_15_20_q  $ (!Xd_0__inst_mult_15_21_q )))))

	.dataa(!Xd_0__inst_mult_15_20_q ),
	.datab(!Xd_0__inst_mult_15_21_q ),
	.datac(!Xd_0__inst_mult_15_22_q ),
	.datad(!Xd_0__inst_mult_15_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_233 ),
	.sharein(Xd_0__inst_mult_15_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_236 ),
	.cout(Xd_0__inst_mult_15_237 ),
	.shareout(Xd_0__inst_mult_15_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_76 (
// Equation(s):
// Xd_0__inst_mult_10_216  = SUM(( !Xd_0__inst_mult_10_20_q  $ (!Xd_0__inst_mult_10_21_q  $ (((Xd_0__inst_mult_10_22_q  & Xd_0__inst_mult_10_23_q )))) ) + ( Xd_0__inst_mult_10_214  ) + ( Xd_0__inst_mult_10_213  ))
// Xd_0__inst_mult_10_217  = CARRY(( !Xd_0__inst_mult_10_20_q  $ (!Xd_0__inst_mult_10_21_q  $ (((Xd_0__inst_mult_10_22_q  & Xd_0__inst_mult_10_23_q )))) ) + ( Xd_0__inst_mult_10_214  ) + ( Xd_0__inst_mult_10_213  ))
// Xd_0__inst_mult_10_218  = SHARE((Xd_0__inst_mult_10_22_q  & (Xd_0__inst_mult_10_23_q  & (!Xd_0__inst_mult_10_20_q  $ (!Xd_0__inst_mult_10_21_q )))))

	.dataa(!Xd_0__inst_mult_10_20_q ),
	.datab(!Xd_0__inst_mult_10_21_q ),
	.datac(!Xd_0__inst_mult_10_22_q ),
	.datad(!Xd_0__inst_mult_10_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_213 ),
	.sharein(Xd_0__inst_mult_10_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_216 ),
	.cout(Xd_0__inst_mult_10_217 ),
	.shareout(Xd_0__inst_mult_10_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_80 (
// Equation(s):
// Xd_0__inst_mult_11_220  = SUM(( !Xd_0__inst_mult_11_20_q  $ (!Xd_0__inst_mult_11_21_q  $ (((Xd_0__inst_mult_11_22_q  & Xd_0__inst_mult_11_23_q )))) ) + ( Xd_0__inst_mult_11_218  ) + ( Xd_0__inst_mult_11_217  ))
// Xd_0__inst_mult_11_221  = CARRY(( !Xd_0__inst_mult_11_20_q  $ (!Xd_0__inst_mult_11_21_q  $ (((Xd_0__inst_mult_11_22_q  & Xd_0__inst_mult_11_23_q )))) ) + ( Xd_0__inst_mult_11_218  ) + ( Xd_0__inst_mult_11_217  ))
// Xd_0__inst_mult_11_222  = SHARE((Xd_0__inst_mult_11_22_q  & (Xd_0__inst_mult_11_23_q  & (!Xd_0__inst_mult_11_20_q  $ (!Xd_0__inst_mult_11_21_q )))))

	.dataa(!Xd_0__inst_mult_11_20_q ),
	.datab(!Xd_0__inst_mult_11_21_q ),
	.datac(!Xd_0__inst_mult_11_22_q ),
	.datad(!Xd_0__inst_mult_11_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_217 ),
	.sharein(Xd_0__inst_mult_11_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_220 ),
	.cout(Xd_0__inst_mult_11_221 ),
	.shareout(Xd_0__inst_mult_11_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_80 (
// Equation(s):
// Xd_0__inst_mult_8_220  = SUM(( !Xd_0__inst_mult_8_20_q  $ (!Xd_0__inst_mult_8_21_q  $ (((Xd_0__inst_mult_8_22_q  & Xd_0__inst_mult_8_23_q )))) ) + ( Xd_0__inst_mult_8_218  ) + ( Xd_0__inst_mult_8_217  ))
// Xd_0__inst_mult_8_221  = CARRY(( !Xd_0__inst_mult_8_20_q  $ (!Xd_0__inst_mult_8_21_q  $ (((Xd_0__inst_mult_8_22_q  & Xd_0__inst_mult_8_23_q )))) ) + ( Xd_0__inst_mult_8_218  ) + ( Xd_0__inst_mult_8_217  ))
// Xd_0__inst_mult_8_222  = SHARE((Xd_0__inst_mult_8_22_q  & (Xd_0__inst_mult_8_23_q  & (!Xd_0__inst_mult_8_20_q  $ (!Xd_0__inst_mult_8_21_q )))))

	.dataa(!Xd_0__inst_mult_8_20_q ),
	.datab(!Xd_0__inst_mult_8_21_q ),
	.datac(!Xd_0__inst_mult_8_22_q ),
	.datad(!Xd_0__inst_mult_8_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_217 ),
	.sharein(Xd_0__inst_mult_8_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_220 ),
	.cout(Xd_0__inst_mult_8_221 ),
	.shareout(Xd_0__inst_mult_8_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_76 (
// Equation(s):
// Xd_0__inst_mult_9_216  = SUM(( !Xd_0__inst_mult_9_20_q  $ (!Xd_0__inst_mult_9_21_q  $ (((Xd_0__inst_mult_9_22_q  & Xd_0__inst_mult_9_23_q )))) ) + ( Xd_0__inst_mult_9_214  ) + ( Xd_0__inst_mult_9_213  ))
// Xd_0__inst_mult_9_217  = CARRY(( !Xd_0__inst_mult_9_20_q  $ (!Xd_0__inst_mult_9_21_q  $ (((Xd_0__inst_mult_9_22_q  & Xd_0__inst_mult_9_23_q )))) ) + ( Xd_0__inst_mult_9_214  ) + ( Xd_0__inst_mult_9_213  ))
// Xd_0__inst_mult_9_218  = SHARE((Xd_0__inst_mult_9_22_q  & (Xd_0__inst_mult_9_23_q  & (!Xd_0__inst_mult_9_20_q  $ (!Xd_0__inst_mult_9_21_q )))))

	.dataa(!Xd_0__inst_mult_9_20_q ),
	.datab(!Xd_0__inst_mult_9_21_q ),
	.datac(!Xd_0__inst_mult_9_22_q ),
	.datad(!Xd_0__inst_mult_9_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_213 ),
	.sharein(Xd_0__inst_mult_9_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_216 ),
	.cout(Xd_0__inst_mult_9_217 ),
	.shareout(Xd_0__inst_mult_9_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_76 (
// Equation(s):
// Xd_0__inst_mult_6_216  = SUM(( !Xd_0__inst_mult_6_20_q  $ (!Xd_0__inst_mult_6_21_q  $ (((Xd_0__inst_mult_6_22_q  & Xd_0__inst_mult_6_23_q )))) ) + ( Xd_0__inst_mult_6_214  ) + ( Xd_0__inst_mult_6_213  ))
// Xd_0__inst_mult_6_217  = CARRY(( !Xd_0__inst_mult_6_20_q  $ (!Xd_0__inst_mult_6_21_q  $ (((Xd_0__inst_mult_6_22_q  & Xd_0__inst_mult_6_23_q )))) ) + ( Xd_0__inst_mult_6_214  ) + ( Xd_0__inst_mult_6_213  ))
// Xd_0__inst_mult_6_218  = SHARE((Xd_0__inst_mult_6_22_q  & (Xd_0__inst_mult_6_23_q  & (!Xd_0__inst_mult_6_20_q  $ (!Xd_0__inst_mult_6_21_q )))))

	.dataa(!Xd_0__inst_mult_6_20_q ),
	.datab(!Xd_0__inst_mult_6_21_q ),
	.datac(!Xd_0__inst_mult_6_22_q ),
	.datad(!Xd_0__inst_mult_6_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_213 ),
	.sharein(Xd_0__inst_mult_6_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_216 ),
	.cout(Xd_0__inst_mult_6_217 ),
	.shareout(Xd_0__inst_mult_6_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_74 (
// Equation(s):
// Xd_0__inst_mult_7_208  = SUM(( !Xd_0__inst_mult_7_20_q  $ (!Xd_0__inst_mult_7_21_q  $ (((Xd_0__inst_mult_7_22_q  & Xd_0__inst_mult_7_23_q )))) ) + ( Xd_0__inst_mult_7_206  ) + ( Xd_0__inst_mult_7_205  ))
// Xd_0__inst_mult_7_209  = CARRY(( !Xd_0__inst_mult_7_20_q  $ (!Xd_0__inst_mult_7_21_q  $ (((Xd_0__inst_mult_7_22_q  & Xd_0__inst_mult_7_23_q )))) ) + ( Xd_0__inst_mult_7_206  ) + ( Xd_0__inst_mult_7_205  ))
// Xd_0__inst_mult_7_210  = SHARE((Xd_0__inst_mult_7_22_q  & (Xd_0__inst_mult_7_23_q  & (!Xd_0__inst_mult_7_20_q  $ (!Xd_0__inst_mult_7_21_q )))))

	.dataa(!Xd_0__inst_mult_7_20_q ),
	.datab(!Xd_0__inst_mult_7_21_q ),
	.datac(!Xd_0__inst_mult_7_22_q ),
	.datad(!Xd_0__inst_mult_7_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_205 ),
	.sharein(Xd_0__inst_mult_7_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_208 ),
	.cout(Xd_0__inst_mult_7_209 ),
	.shareout(Xd_0__inst_mult_7_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_84 (
// Equation(s):
// Xd_0__inst_mult_4_236  = SUM(( !Xd_0__inst_mult_4_20_q  $ (!Xd_0__inst_mult_4_21_q  $ (((Xd_0__inst_mult_4_22_q  & Xd_0__inst_mult_4_23_q )))) ) + ( Xd_0__inst_mult_4_234  ) + ( Xd_0__inst_mult_4_233  ))
// Xd_0__inst_mult_4_237  = CARRY(( !Xd_0__inst_mult_4_20_q  $ (!Xd_0__inst_mult_4_21_q  $ (((Xd_0__inst_mult_4_22_q  & Xd_0__inst_mult_4_23_q )))) ) + ( Xd_0__inst_mult_4_234  ) + ( Xd_0__inst_mult_4_233  ))
// Xd_0__inst_mult_4_238  = SHARE((Xd_0__inst_mult_4_22_q  & (Xd_0__inst_mult_4_23_q  & (!Xd_0__inst_mult_4_20_q  $ (!Xd_0__inst_mult_4_21_q )))))

	.dataa(!Xd_0__inst_mult_4_20_q ),
	.datab(!Xd_0__inst_mult_4_21_q ),
	.datac(!Xd_0__inst_mult_4_22_q ),
	.datad(!Xd_0__inst_mult_4_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_233 ),
	.sharein(Xd_0__inst_mult_4_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_236 ),
	.cout(Xd_0__inst_mult_4_237 ),
	.shareout(Xd_0__inst_mult_4_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_74 (
// Equation(s):
// Xd_0__inst_mult_5_208  = SUM(( !Xd_0__inst_mult_5_20_q  $ (!Xd_0__inst_mult_5_21_q  $ (((Xd_0__inst_mult_5_22_q  & Xd_0__inst_mult_5_23_q )))) ) + ( Xd_0__inst_mult_5_206  ) + ( Xd_0__inst_mult_5_205  ))
// Xd_0__inst_mult_5_209  = CARRY(( !Xd_0__inst_mult_5_20_q  $ (!Xd_0__inst_mult_5_21_q  $ (((Xd_0__inst_mult_5_22_q  & Xd_0__inst_mult_5_23_q )))) ) + ( Xd_0__inst_mult_5_206  ) + ( Xd_0__inst_mult_5_205  ))
// Xd_0__inst_mult_5_210  = SHARE((Xd_0__inst_mult_5_22_q  & (Xd_0__inst_mult_5_23_q  & (!Xd_0__inst_mult_5_20_q  $ (!Xd_0__inst_mult_5_21_q )))))

	.dataa(!Xd_0__inst_mult_5_20_q ),
	.datab(!Xd_0__inst_mult_5_21_q ),
	.datac(!Xd_0__inst_mult_5_22_q ),
	.datad(!Xd_0__inst_mult_5_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_205 ),
	.sharein(Xd_0__inst_mult_5_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_208 ),
	.cout(Xd_0__inst_mult_5_209 ),
	.shareout(Xd_0__inst_mult_5_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_78 (
// Equation(s):
// Xd_0__inst_mult_2_212  = SUM(( !Xd_0__inst_mult_2_20_q  $ (!Xd_0__inst_mult_2_21_q  $ (((Xd_0__inst_mult_2_22_q  & Xd_0__inst_mult_2_23_q )))) ) + ( Xd_0__inst_mult_2_210  ) + ( Xd_0__inst_mult_2_209  ))
// Xd_0__inst_mult_2_213  = CARRY(( !Xd_0__inst_mult_2_20_q  $ (!Xd_0__inst_mult_2_21_q  $ (((Xd_0__inst_mult_2_22_q  & Xd_0__inst_mult_2_23_q )))) ) + ( Xd_0__inst_mult_2_210  ) + ( Xd_0__inst_mult_2_209  ))
// Xd_0__inst_mult_2_214  = SHARE((Xd_0__inst_mult_2_22_q  & (Xd_0__inst_mult_2_23_q  & (!Xd_0__inst_mult_2_20_q  $ (!Xd_0__inst_mult_2_21_q )))))

	.dataa(!Xd_0__inst_mult_2_20_q ),
	.datab(!Xd_0__inst_mult_2_21_q ),
	.datac(!Xd_0__inst_mult_2_22_q ),
	.datad(!Xd_0__inst_mult_2_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_209 ),
	.sharein(Xd_0__inst_mult_2_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_212 ),
	.cout(Xd_0__inst_mult_2_213 ),
	.shareout(Xd_0__inst_mult_2_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_74 (
// Equation(s):
// Xd_0__inst_mult_3_208  = SUM(( !Xd_0__inst_mult_3_20_q  $ (!Xd_0__inst_mult_3_21_q  $ (((Xd_0__inst_mult_3_22_q  & Xd_0__inst_mult_3_23_q )))) ) + ( Xd_0__inst_mult_3_206  ) + ( Xd_0__inst_mult_3_205  ))
// Xd_0__inst_mult_3_209  = CARRY(( !Xd_0__inst_mult_3_20_q  $ (!Xd_0__inst_mult_3_21_q  $ (((Xd_0__inst_mult_3_22_q  & Xd_0__inst_mult_3_23_q )))) ) + ( Xd_0__inst_mult_3_206  ) + ( Xd_0__inst_mult_3_205  ))
// Xd_0__inst_mult_3_210  = SHARE((Xd_0__inst_mult_3_22_q  & (Xd_0__inst_mult_3_23_q  & (!Xd_0__inst_mult_3_20_q  $ (!Xd_0__inst_mult_3_21_q )))))

	.dataa(!Xd_0__inst_mult_3_20_q ),
	.datab(!Xd_0__inst_mult_3_21_q ),
	.datac(!Xd_0__inst_mult_3_22_q ),
	.datad(!Xd_0__inst_mult_3_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_205 ),
	.sharein(Xd_0__inst_mult_3_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_208 ),
	.cout(Xd_0__inst_mult_3_209 ),
	.shareout(Xd_0__inst_mult_3_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_78 (
// Equation(s):
// Xd_0__inst_mult_0_212  = SUM(( !Xd_0__inst_mult_0_20_q  $ (!Xd_0__inst_mult_0_21_q  $ (((Xd_0__inst_mult_0_22_q  & Xd_0__inst_mult_0_23_q )))) ) + ( Xd_0__inst_mult_0_210  ) + ( Xd_0__inst_mult_0_209  ))
// Xd_0__inst_mult_0_213  = CARRY(( !Xd_0__inst_mult_0_20_q  $ (!Xd_0__inst_mult_0_21_q  $ (((Xd_0__inst_mult_0_22_q  & Xd_0__inst_mult_0_23_q )))) ) + ( Xd_0__inst_mult_0_210  ) + ( Xd_0__inst_mult_0_209  ))
// Xd_0__inst_mult_0_214  = SHARE((Xd_0__inst_mult_0_22_q  & (Xd_0__inst_mult_0_23_q  & (!Xd_0__inst_mult_0_20_q  $ (!Xd_0__inst_mult_0_21_q )))))

	.dataa(!Xd_0__inst_mult_0_20_q ),
	.datab(!Xd_0__inst_mult_0_21_q ),
	.datac(!Xd_0__inst_mult_0_22_q ),
	.datad(!Xd_0__inst_mult_0_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_209 ),
	.sharein(Xd_0__inst_mult_0_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_212 ),
	.cout(Xd_0__inst_mult_0_213 ),
	.shareout(Xd_0__inst_mult_0_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_78 (
// Equation(s):
// Xd_0__inst_mult_1_212  = SUM(( !Xd_0__inst_mult_1_20_q  $ (!Xd_0__inst_mult_1_21_q  $ (((Xd_0__inst_mult_1_22_q  & Xd_0__inst_mult_1_23_q )))) ) + ( Xd_0__inst_mult_1_210  ) + ( Xd_0__inst_mult_1_209  ))
// Xd_0__inst_mult_1_213  = CARRY(( !Xd_0__inst_mult_1_20_q  $ (!Xd_0__inst_mult_1_21_q  $ (((Xd_0__inst_mult_1_22_q  & Xd_0__inst_mult_1_23_q )))) ) + ( Xd_0__inst_mult_1_210  ) + ( Xd_0__inst_mult_1_209  ))
// Xd_0__inst_mult_1_214  = SHARE((Xd_0__inst_mult_1_22_q  & (Xd_0__inst_mult_1_23_q  & (!Xd_0__inst_mult_1_20_q  $ (!Xd_0__inst_mult_1_21_q )))))

	.dataa(!Xd_0__inst_mult_1_20_q ),
	.datab(!Xd_0__inst_mult_1_21_q ),
	.datac(!Xd_0__inst_mult_1_22_q ),
	.datad(!Xd_0__inst_mult_1_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_209 ),
	.sharein(Xd_0__inst_mult_1_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_212 ),
	.cout(Xd_0__inst_mult_1_213 ),
	.shareout(Xd_0__inst_mult_1_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_81 (
// Equation(s):
// Xd_0__inst_mult_12_236  = SUM(( !Xd_0__inst_mult_12_24_q  $ (!Xd_0__inst_mult_12_25_q  $ (((Xd_0__inst_mult_12_20_q  & Xd_0__inst_mult_12_21_q )))) ) + ( Xd_0__inst_mult_12_234  ) + ( Xd_0__inst_mult_12_233  ))
// Xd_0__inst_mult_12_237  = CARRY(( !Xd_0__inst_mult_12_24_q  $ (!Xd_0__inst_mult_12_25_q  $ (((Xd_0__inst_mult_12_20_q  & Xd_0__inst_mult_12_21_q )))) ) + ( Xd_0__inst_mult_12_234  ) + ( Xd_0__inst_mult_12_233  ))
// Xd_0__inst_mult_12_238  = SHARE((Xd_0__inst_mult_12_20_q  & (Xd_0__inst_mult_12_21_q  & (!Xd_0__inst_mult_12_24_q  $ (!Xd_0__inst_mult_12_25_q )))))

	.dataa(!Xd_0__inst_mult_12_24_q ),
	.datab(!Xd_0__inst_mult_12_25_q ),
	.datac(!Xd_0__inst_mult_12_20_q ),
	.datad(!Xd_0__inst_mult_12_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_233 ),
	.sharein(Xd_0__inst_mult_12_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_236 ),
	.cout(Xd_0__inst_mult_12_237 ),
	.shareout(Xd_0__inst_mult_12_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_81 (
// Equation(s):
// Xd_0__inst_mult_13_224  = SUM(( !Xd_0__inst_mult_13_24_q  $ (!Xd_0__inst_mult_13_25_q  $ (((Xd_0__inst_mult_13_20_q  & Xd_0__inst_mult_13_21_q )))) ) + ( Xd_0__inst_mult_13_222  ) + ( Xd_0__inst_mult_13_221  ))
// Xd_0__inst_mult_13_225  = CARRY(( !Xd_0__inst_mult_13_24_q  $ (!Xd_0__inst_mult_13_25_q  $ (((Xd_0__inst_mult_13_20_q  & Xd_0__inst_mult_13_21_q )))) ) + ( Xd_0__inst_mult_13_222  ) + ( Xd_0__inst_mult_13_221  ))
// Xd_0__inst_mult_13_226  = SHARE((Xd_0__inst_mult_13_20_q  & (Xd_0__inst_mult_13_21_q  & (!Xd_0__inst_mult_13_24_q  $ (!Xd_0__inst_mult_13_25_q )))))

	.dataa(!Xd_0__inst_mult_13_24_q ),
	.datab(!Xd_0__inst_mult_13_25_q ),
	.datac(!Xd_0__inst_mult_13_20_q ),
	.datad(!Xd_0__inst_mult_13_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_221 ),
	.sharein(Xd_0__inst_mult_13_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_224 ),
	.cout(Xd_0__inst_mult_13_225 ),
	.shareout(Xd_0__inst_mult_13_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_85 (
// Equation(s):
// Xd_0__inst_mult_14_240  = SUM(( !Xd_0__inst_mult_14_24_q  $ (!Xd_0__inst_mult_14_25_q  $ (((Xd_0__inst_mult_14_20_q  & Xd_0__inst_mult_14_21_q )))) ) + ( Xd_0__inst_mult_14_238  ) + ( Xd_0__inst_mult_14_237  ))
// Xd_0__inst_mult_14_241  = CARRY(( !Xd_0__inst_mult_14_24_q  $ (!Xd_0__inst_mult_14_25_q  $ (((Xd_0__inst_mult_14_20_q  & Xd_0__inst_mult_14_21_q )))) ) + ( Xd_0__inst_mult_14_238  ) + ( Xd_0__inst_mult_14_237  ))
// Xd_0__inst_mult_14_242  = SHARE((Xd_0__inst_mult_14_20_q  & (Xd_0__inst_mult_14_21_q  & (!Xd_0__inst_mult_14_24_q  $ (!Xd_0__inst_mult_14_25_q )))))

	.dataa(!Xd_0__inst_mult_14_24_q ),
	.datab(!Xd_0__inst_mult_14_25_q ),
	.datac(!Xd_0__inst_mult_14_20_q ),
	.datad(!Xd_0__inst_mult_14_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_237 ),
	.sharein(Xd_0__inst_mult_14_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_240 ),
	.cout(Xd_0__inst_mult_14_241 ),
	.shareout(Xd_0__inst_mult_14_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_85 (
// Equation(s):
// Xd_0__inst_mult_15_240  = SUM(( !Xd_0__inst_mult_15_24_q  $ (!Xd_0__inst_mult_15_25_q  $ (((Xd_0__inst_mult_15_20_q  & Xd_0__inst_mult_15_21_q )))) ) + ( Xd_0__inst_mult_15_238  ) + ( Xd_0__inst_mult_15_237  ))
// Xd_0__inst_mult_15_241  = CARRY(( !Xd_0__inst_mult_15_24_q  $ (!Xd_0__inst_mult_15_25_q  $ (((Xd_0__inst_mult_15_20_q  & Xd_0__inst_mult_15_21_q )))) ) + ( Xd_0__inst_mult_15_238  ) + ( Xd_0__inst_mult_15_237  ))
// Xd_0__inst_mult_15_242  = SHARE((Xd_0__inst_mult_15_20_q  & (Xd_0__inst_mult_15_21_q  & (!Xd_0__inst_mult_15_24_q  $ (!Xd_0__inst_mult_15_25_q )))))

	.dataa(!Xd_0__inst_mult_15_24_q ),
	.datab(!Xd_0__inst_mult_15_25_q ),
	.datac(!Xd_0__inst_mult_15_20_q ),
	.datad(!Xd_0__inst_mult_15_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_237 ),
	.sharein(Xd_0__inst_mult_15_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_240 ),
	.cout(Xd_0__inst_mult_15_241 ),
	.shareout(Xd_0__inst_mult_15_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_77 (
// Equation(s):
// Xd_0__inst_mult_10_220  = SUM(( !Xd_0__inst_mult_10_24_q  $ (!Xd_0__inst_mult_10_25_q  $ (((Xd_0__inst_mult_10_20_q  & Xd_0__inst_mult_10_21_q )))) ) + ( Xd_0__inst_mult_10_218  ) + ( Xd_0__inst_mult_10_217  ))
// Xd_0__inst_mult_10_221  = CARRY(( !Xd_0__inst_mult_10_24_q  $ (!Xd_0__inst_mult_10_25_q  $ (((Xd_0__inst_mult_10_20_q  & Xd_0__inst_mult_10_21_q )))) ) + ( Xd_0__inst_mult_10_218  ) + ( Xd_0__inst_mult_10_217  ))
// Xd_0__inst_mult_10_222  = SHARE((Xd_0__inst_mult_10_20_q  & (Xd_0__inst_mult_10_21_q  & (!Xd_0__inst_mult_10_24_q  $ (!Xd_0__inst_mult_10_25_q )))))

	.dataa(!Xd_0__inst_mult_10_24_q ),
	.datab(!Xd_0__inst_mult_10_25_q ),
	.datac(!Xd_0__inst_mult_10_20_q ),
	.datad(!Xd_0__inst_mult_10_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_217 ),
	.sharein(Xd_0__inst_mult_10_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_220 ),
	.cout(Xd_0__inst_mult_10_221 ),
	.shareout(Xd_0__inst_mult_10_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_81 (
// Equation(s):
// Xd_0__inst_mult_11_224  = SUM(( !Xd_0__inst_mult_11_24_q  $ (!Xd_0__inst_mult_11_25_q  $ (((Xd_0__inst_mult_11_20_q  & Xd_0__inst_mult_11_21_q )))) ) + ( Xd_0__inst_mult_11_222  ) + ( Xd_0__inst_mult_11_221  ))
// Xd_0__inst_mult_11_225  = CARRY(( !Xd_0__inst_mult_11_24_q  $ (!Xd_0__inst_mult_11_25_q  $ (((Xd_0__inst_mult_11_20_q  & Xd_0__inst_mult_11_21_q )))) ) + ( Xd_0__inst_mult_11_222  ) + ( Xd_0__inst_mult_11_221  ))
// Xd_0__inst_mult_11_226  = SHARE((Xd_0__inst_mult_11_20_q  & (Xd_0__inst_mult_11_21_q  & (!Xd_0__inst_mult_11_24_q  $ (!Xd_0__inst_mult_11_25_q )))))

	.dataa(!Xd_0__inst_mult_11_24_q ),
	.datab(!Xd_0__inst_mult_11_25_q ),
	.datac(!Xd_0__inst_mult_11_20_q ),
	.datad(!Xd_0__inst_mult_11_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_221 ),
	.sharein(Xd_0__inst_mult_11_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_224 ),
	.cout(Xd_0__inst_mult_11_225 ),
	.shareout(Xd_0__inst_mult_11_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_81 (
// Equation(s):
// Xd_0__inst_mult_8_224  = SUM(( !Xd_0__inst_mult_8_24_q  $ (!Xd_0__inst_mult_8_25_q  $ (((Xd_0__inst_mult_8_20_q  & Xd_0__inst_mult_8_21_q )))) ) + ( Xd_0__inst_mult_8_222  ) + ( Xd_0__inst_mult_8_221  ))
// Xd_0__inst_mult_8_225  = CARRY(( !Xd_0__inst_mult_8_24_q  $ (!Xd_0__inst_mult_8_25_q  $ (((Xd_0__inst_mult_8_20_q  & Xd_0__inst_mult_8_21_q )))) ) + ( Xd_0__inst_mult_8_222  ) + ( Xd_0__inst_mult_8_221  ))
// Xd_0__inst_mult_8_226  = SHARE((Xd_0__inst_mult_8_20_q  & (Xd_0__inst_mult_8_21_q  & (!Xd_0__inst_mult_8_24_q  $ (!Xd_0__inst_mult_8_25_q )))))

	.dataa(!Xd_0__inst_mult_8_24_q ),
	.datab(!Xd_0__inst_mult_8_25_q ),
	.datac(!Xd_0__inst_mult_8_20_q ),
	.datad(!Xd_0__inst_mult_8_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_221 ),
	.sharein(Xd_0__inst_mult_8_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_224 ),
	.cout(Xd_0__inst_mult_8_225 ),
	.shareout(Xd_0__inst_mult_8_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_77 (
// Equation(s):
// Xd_0__inst_mult_9_220  = SUM(( !Xd_0__inst_mult_9_24_q  $ (!Xd_0__inst_mult_9_25_q  $ (((Xd_0__inst_mult_9_20_q  & Xd_0__inst_mult_9_21_q )))) ) + ( Xd_0__inst_mult_9_218  ) + ( Xd_0__inst_mult_9_217  ))
// Xd_0__inst_mult_9_221  = CARRY(( !Xd_0__inst_mult_9_24_q  $ (!Xd_0__inst_mult_9_25_q  $ (((Xd_0__inst_mult_9_20_q  & Xd_0__inst_mult_9_21_q )))) ) + ( Xd_0__inst_mult_9_218  ) + ( Xd_0__inst_mult_9_217  ))
// Xd_0__inst_mult_9_222  = SHARE((Xd_0__inst_mult_9_20_q  & (Xd_0__inst_mult_9_21_q  & (!Xd_0__inst_mult_9_24_q  $ (!Xd_0__inst_mult_9_25_q )))))

	.dataa(!Xd_0__inst_mult_9_24_q ),
	.datab(!Xd_0__inst_mult_9_25_q ),
	.datac(!Xd_0__inst_mult_9_20_q ),
	.datad(!Xd_0__inst_mult_9_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_217 ),
	.sharein(Xd_0__inst_mult_9_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_220 ),
	.cout(Xd_0__inst_mult_9_221 ),
	.shareout(Xd_0__inst_mult_9_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_77 (
// Equation(s):
// Xd_0__inst_mult_6_220  = SUM(( !Xd_0__inst_mult_6_24_q  $ (!Xd_0__inst_mult_6_25_q  $ (((Xd_0__inst_mult_6_20_q  & Xd_0__inst_mult_6_21_q )))) ) + ( Xd_0__inst_mult_6_218  ) + ( Xd_0__inst_mult_6_217  ))
// Xd_0__inst_mult_6_221  = CARRY(( !Xd_0__inst_mult_6_24_q  $ (!Xd_0__inst_mult_6_25_q  $ (((Xd_0__inst_mult_6_20_q  & Xd_0__inst_mult_6_21_q )))) ) + ( Xd_0__inst_mult_6_218  ) + ( Xd_0__inst_mult_6_217  ))
// Xd_0__inst_mult_6_222  = SHARE((Xd_0__inst_mult_6_20_q  & (Xd_0__inst_mult_6_21_q  & (!Xd_0__inst_mult_6_24_q  $ (!Xd_0__inst_mult_6_25_q )))))

	.dataa(!Xd_0__inst_mult_6_24_q ),
	.datab(!Xd_0__inst_mult_6_25_q ),
	.datac(!Xd_0__inst_mult_6_20_q ),
	.datad(!Xd_0__inst_mult_6_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_217 ),
	.sharein(Xd_0__inst_mult_6_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_220 ),
	.cout(Xd_0__inst_mult_6_221 ),
	.shareout(Xd_0__inst_mult_6_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_75 (
// Equation(s):
// Xd_0__inst_mult_7_212  = SUM(( !Xd_0__inst_mult_7_24_q  $ (!Xd_0__inst_mult_7_25_q  $ (((Xd_0__inst_mult_7_20_q  & Xd_0__inst_mult_7_21_q )))) ) + ( Xd_0__inst_mult_7_210  ) + ( Xd_0__inst_mult_7_209  ))
// Xd_0__inst_mult_7_213  = CARRY(( !Xd_0__inst_mult_7_24_q  $ (!Xd_0__inst_mult_7_25_q  $ (((Xd_0__inst_mult_7_20_q  & Xd_0__inst_mult_7_21_q )))) ) + ( Xd_0__inst_mult_7_210  ) + ( Xd_0__inst_mult_7_209  ))
// Xd_0__inst_mult_7_214  = SHARE((Xd_0__inst_mult_7_20_q  & (Xd_0__inst_mult_7_21_q  & (!Xd_0__inst_mult_7_24_q  $ (!Xd_0__inst_mult_7_25_q )))))

	.dataa(!Xd_0__inst_mult_7_24_q ),
	.datab(!Xd_0__inst_mult_7_25_q ),
	.datac(!Xd_0__inst_mult_7_20_q ),
	.datad(!Xd_0__inst_mult_7_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_209 ),
	.sharein(Xd_0__inst_mult_7_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_212 ),
	.cout(Xd_0__inst_mult_7_213 ),
	.shareout(Xd_0__inst_mult_7_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_85 (
// Equation(s):
// Xd_0__inst_mult_4_240  = SUM(( !Xd_0__inst_mult_4_24_q  $ (!Xd_0__inst_mult_4_25_q  $ (((Xd_0__inst_mult_4_20_q  & Xd_0__inst_mult_4_21_q )))) ) + ( Xd_0__inst_mult_4_238  ) + ( Xd_0__inst_mult_4_237  ))
// Xd_0__inst_mult_4_241  = CARRY(( !Xd_0__inst_mult_4_24_q  $ (!Xd_0__inst_mult_4_25_q  $ (((Xd_0__inst_mult_4_20_q  & Xd_0__inst_mult_4_21_q )))) ) + ( Xd_0__inst_mult_4_238  ) + ( Xd_0__inst_mult_4_237  ))
// Xd_0__inst_mult_4_242  = SHARE((Xd_0__inst_mult_4_20_q  & (Xd_0__inst_mult_4_21_q  & (!Xd_0__inst_mult_4_24_q  $ (!Xd_0__inst_mult_4_25_q )))))

	.dataa(!Xd_0__inst_mult_4_24_q ),
	.datab(!Xd_0__inst_mult_4_25_q ),
	.datac(!Xd_0__inst_mult_4_20_q ),
	.datad(!Xd_0__inst_mult_4_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_237 ),
	.sharein(Xd_0__inst_mult_4_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_240 ),
	.cout(Xd_0__inst_mult_4_241 ),
	.shareout(Xd_0__inst_mult_4_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_75 (
// Equation(s):
// Xd_0__inst_mult_5_212  = SUM(( !Xd_0__inst_mult_5_24_q  $ (!Xd_0__inst_mult_5_25_q  $ (((Xd_0__inst_mult_5_20_q  & Xd_0__inst_mult_5_21_q )))) ) + ( Xd_0__inst_mult_5_210  ) + ( Xd_0__inst_mult_5_209  ))
// Xd_0__inst_mult_5_213  = CARRY(( !Xd_0__inst_mult_5_24_q  $ (!Xd_0__inst_mult_5_25_q  $ (((Xd_0__inst_mult_5_20_q  & Xd_0__inst_mult_5_21_q )))) ) + ( Xd_0__inst_mult_5_210  ) + ( Xd_0__inst_mult_5_209  ))
// Xd_0__inst_mult_5_214  = SHARE((Xd_0__inst_mult_5_20_q  & (Xd_0__inst_mult_5_21_q  & (!Xd_0__inst_mult_5_24_q  $ (!Xd_0__inst_mult_5_25_q )))))

	.dataa(!Xd_0__inst_mult_5_24_q ),
	.datab(!Xd_0__inst_mult_5_25_q ),
	.datac(!Xd_0__inst_mult_5_20_q ),
	.datad(!Xd_0__inst_mult_5_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_209 ),
	.sharein(Xd_0__inst_mult_5_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_212 ),
	.cout(Xd_0__inst_mult_5_213 ),
	.shareout(Xd_0__inst_mult_5_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_79 (
// Equation(s):
// Xd_0__inst_mult_2_216  = SUM(( !Xd_0__inst_mult_2_24_q  $ (!Xd_0__inst_mult_2_25_q  $ (((Xd_0__inst_mult_2_20_q  & Xd_0__inst_mult_2_21_q )))) ) + ( Xd_0__inst_mult_2_214  ) + ( Xd_0__inst_mult_2_213  ))
// Xd_0__inst_mult_2_217  = CARRY(( !Xd_0__inst_mult_2_24_q  $ (!Xd_0__inst_mult_2_25_q  $ (((Xd_0__inst_mult_2_20_q  & Xd_0__inst_mult_2_21_q )))) ) + ( Xd_0__inst_mult_2_214  ) + ( Xd_0__inst_mult_2_213  ))
// Xd_0__inst_mult_2_218  = SHARE((Xd_0__inst_mult_2_20_q  & (Xd_0__inst_mult_2_21_q  & (!Xd_0__inst_mult_2_24_q  $ (!Xd_0__inst_mult_2_25_q )))))

	.dataa(!Xd_0__inst_mult_2_24_q ),
	.datab(!Xd_0__inst_mult_2_25_q ),
	.datac(!Xd_0__inst_mult_2_20_q ),
	.datad(!Xd_0__inst_mult_2_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_213 ),
	.sharein(Xd_0__inst_mult_2_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_216 ),
	.cout(Xd_0__inst_mult_2_217 ),
	.shareout(Xd_0__inst_mult_2_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_75 (
// Equation(s):
// Xd_0__inst_mult_3_212  = SUM(( !Xd_0__inst_mult_3_24_q  $ (!Xd_0__inst_mult_3_25_q  $ (((Xd_0__inst_mult_3_20_q  & Xd_0__inst_mult_3_21_q )))) ) + ( Xd_0__inst_mult_3_210  ) + ( Xd_0__inst_mult_3_209  ))
// Xd_0__inst_mult_3_213  = CARRY(( !Xd_0__inst_mult_3_24_q  $ (!Xd_0__inst_mult_3_25_q  $ (((Xd_0__inst_mult_3_20_q  & Xd_0__inst_mult_3_21_q )))) ) + ( Xd_0__inst_mult_3_210  ) + ( Xd_0__inst_mult_3_209  ))
// Xd_0__inst_mult_3_214  = SHARE((Xd_0__inst_mult_3_20_q  & (Xd_0__inst_mult_3_21_q  & (!Xd_0__inst_mult_3_24_q  $ (!Xd_0__inst_mult_3_25_q )))))

	.dataa(!Xd_0__inst_mult_3_24_q ),
	.datab(!Xd_0__inst_mult_3_25_q ),
	.datac(!Xd_0__inst_mult_3_20_q ),
	.datad(!Xd_0__inst_mult_3_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_209 ),
	.sharein(Xd_0__inst_mult_3_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_212 ),
	.cout(Xd_0__inst_mult_3_213 ),
	.shareout(Xd_0__inst_mult_3_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_79 (
// Equation(s):
// Xd_0__inst_mult_0_216  = SUM(( !Xd_0__inst_mult_0_24_q  $ (!Xd_0__inst_mult_0_25_q  $ (((Xd_0__inst_mult_0_20_q  & Xd_0__inst_mult_0_21_q )))) ) + ( Xd_0__inst_mult_0_214  ) + ( Xd_0__inst_mult_0_213  ))
// Xd_0__inst_mult_0_217  = CARRY(( !Xd_0__inst_mult_0_24_q  $ (!Xd_0__inst_mult_0_25_q  $ (((Xd_0__inst_mult_0_20_q  & Xd_0__inst_mult_0_21_q )))) ) + ( Xd_0__inst_mult_0_214  ) + ( Xd_0__inst_mult_0_213  ))
// Xd_0__inst_mult_0_218  = SHARE((Xd_0__inst_mult_0_20_q  & (Xd_0__inst_mult_0_21_q  & (!Xd_0__inst_mult_0_24_q  $ (!Xd_0__inst_mult_0_25_q )))))

	.dataa(!Xd_0__inst_mult_0_24_q ),
	.datab(!Xd_0__inst_mult_0_25_q ),
	.datac(!Xd_0__inst_mult_0_20_q ),
	.datad(!Xd_0__inst_mult_0_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_213 ),
	.sharein(Xd_0__inst_mult_0_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_216 ),
	.cout(Xd_0__inst_mult_0_217 ),
	.shareout(Xd_0__inst_mult_0_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_79 (
// Equation(s):
// Xd_0__inst_mult_1_216  = SUM(( !Xd_0__inst_mult_1_24_q  $ (!Xd_0__inst_mult_1_25_q  $ (((Xd_0__inst_mult_1_20_q  & Xd_0__inst_mult_1_21_q )))) ) + ( Xd_0__inst_mult_1_214  ) + ( Xd_0__inst_mult_1_213  ))
// Xd_0__inst_mult_1_217  = CARRY(( !Xd_0__inst_mult_1_24_q  $ (!Xd_0__inst_mult_1_25_q  $ (((Xd_0__inst_mult_1_20_q  & Xd_0__inst_mult_1_21_q )))) ) + ( Xd_0__inst_mult_1_214  ) + ( Xd_0__inst_mult_1_213  ))
// Xd_0__inst_mult_1_218  = SHARE((Xd_0__inst_mult_1_20_q  & (Xd_0__inst_mult_1_21_q  & (!Xd_0__inst_mult_1_24_q  $ (!Xd_0__inst_mult_1_25_q )))))

	.dataa(!Xd_0__inst_mult_1_24_q ),
	.datab(!Xd_0__inst_mult_1_25_q ),
	.datac(!Xd_0__inst_mult_1_20_q ),
	.datad(!Xd_0__inst_mult_1_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_213 ),
	.sharein(Xd_0__inst_mult_1_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_216 ),
	.cout(Xd_0__inst_mult_1_217 ),
	.shareout(Xd_0__inst_mult_1_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_82 (
// Equation(s):
// Xd_0__inst_mult_12_240  = SUM(( !Xd_0__inst_mult_12_26_q  $ (!Xd_0__inst_mult_12_27_q  $ (((Xd_0__inst_mult_12_24_q  & Xd_0__inst_mult_12_25_q )))) ) + ( Xd_0__inst_mult_12_238  ) + ( Xd_0__inst_mult_12_237  ))
// Xd_0__inst_mult_12_241  = CARRY(( !Xd_0__inst_mult_12_26_q  $ (!Xd_0__inst_mult_12_27_q  $ (((Xd_0__inst_mult_12_24_q  & Xd_0__inst_mult_12_25_q )))) ) + ( Xd_0__inst_mult_12_238  ) + ( Xd_0__inst_mult_12_237  ))
// Xd_0__inst_mult_12_242  = SHARE((Xd_0__inst_mult_12_24_q  & (Xd_0__inst_mult_12_25_q  & (!Xd_0__inst_mult_12_26_q  $ (!Xd_0__inst_mult_12_27_q )))))

	.dataa(!Xd_0__inst_mult_12_26_q ),
	.datab(!Xd_0__inst_mult_12_27_q ),
	.datac(!Xd_0__inst_mult_12_24_q ),
	.datad(!Xd_0__inst_mult_12_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_237 ),
	.sharein(Xd_0__inst_mult_12_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_240 ),
	.cout(Xd_0__inst_mult_12_241 ),
	.shareout(Xd_0__inst_mult_12_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_82 (
// Equation(s):
// Xd_0__inst_mult_13_228  = SUM(( !Xd_0__inst_mult_13_26_q  $ (!Xd_0__inst_mult_13_27_q  $ (((Xd_0__inst_mult_13_24_q  & Xd_0__inst_mult_13_25_q )))) ) + ( Xd_0__inst_mult_13_226  ) + ( Xd_0__inst_mult_13_225  ))
// Xd_0__inst_mult_13_229  = CARRY(( !Xd_0__inst_mult_13_26_q  $ (!Xd_0__inst_mult_13_27_q  $ (((Xd_0__inst_mult_13_24_q  & Xd_0__inst_mult_13_25_q )))) ) + ( Xd_0__inst_mult_13_226  ) + ( Xd_0__inst_mult_13_225  ))
// Xd_0__inst_mult_13_230  = SHARE((Xd_0__inst_mult_13_24_q  & (Xd_0__inst_mult_13_25_q  & (!Xd_0__inst_mult_13_26_q  $ (!Xd_0__inst_mult_13_27_q )))))

	.dataa(!Xd_0__inst_mult_13_26_q ),
	.datab(!Xd_0__inst_mult_13_27_q ),
	.datac(!Xd_0__inst_mult_13_24_q ),
	.datad(!Xd_0__inst_mult_13_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_225 ),
	.sharein(Xd_0__inst_mult_13_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_228 ),
	.cout(Xd_0__inst_mult_13_229 ),
	.shareout(Xd_0__inst_mult_13_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_86 (
// Equation(s):
// Xd_0__inst_mult_14_244  = SUM(( !Xd_0__inst_mult_14_26_q  $ (!Xd_0__inst_mult_14_27_q  $ (((Xd_0__inst_mult_14_24_q  & Xd_0__inst_mult_14_25_q )))) ) + ( Xd_0__inst_mult_14_242  ) + ( Xd_0__inst_mult_14_241  ))
// Xd_0__inst_mult_14_245  = CARRY(( !Xd_0__inst_mult_14_26_q  $ (!Xd_0__inst_mult_14_27_q  $ (((Xd_0__inst_mult_14_24_q  & Xd_0__inst_mult_14_25_q )))) ) + ( Xd_0__inst_mult_14_242  ) + ( Xd_0__inst_mult_14_241  ))
// Xd_0__inst_mult_14_246  = SHARE((Xd_0__inst_mult_14_24_q  & (Xd_0__inst_mult_14_25_q  & (!Xd_0__inst_mult_14_26_q  $ (!Xd_0__inst_mult_14_27_q )))))

	.dataa(!Xd_0__inst_mult_14_26_q ),
	.datab(!Xd_0__inst_mult_14_27_q ),
	.datac(!Xd_0__inst_mult_14_24_q ),
	.datad(!Xd_0__inst_mult_14_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_241 ),
	.sharein(Xd_0__inst_mult_14_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_244 ),
	.cout(Xd_0__inst_mult_14_245 ),
	.shareout(Xd_0__inst_mult_14_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_86 (
// Equation(s):
// Xd_0__inst_mult_15_244  = SUM(( !Xd_0__inst_mult_15_26_q  $ (!Xd_0__inst_mult_15_27_q  $ (((Xd_0__inst_mult_15_24_q  & Xd_0__inst_mult_15_25_q )))) ) + ( Xd_0__inst_mult_15_242  ) + ( Xd_0__inst_mult_15_241  ))
// Xd_0__inst_mult_15_245  = CARRY(( !Xd_0__inst_mult_15_26_q  $ (!Xd_0__inst_mult_15_27_q  $ (((Xd_0__inst_mult_15_24_q  & Xd_0__inst_mult_15_25_q )))) ) + ( Xd_0__inst_mult_15_242  ) + ( Xd_0__inst_mult_15_241  ))
// Xd_0__inst_mult_15_246  = SHARE((Xd_0__inst_mult_15_24_q  & (Xd_0__inst_mult_15_25_q  & (!Xd_0__inst_mult_15_26_q  $ (!Xd_0__inst_mult_15_27_q )))))

	.dataa(!Xd_0__inst_mult_15_26_q ),
	.datab(!Xd_0__inst_mult_15_27_q ),
	.datac(!Xd_0__inst_mult_15_24_q ),
	.datad(!Xd_0__inst_mult_15_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_241 ),
	.sharein(Xd_0__inst_mult_15_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_244 ),
	.cout(Xd_0__inst_mult_15_245 ),
	.shareout(Xd_0__inst_mult_15_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_78 (
// Equation(s):
// Xd_0__inst_mult_10_224  = SUM(( !Xd_0__inst_mult_10_26_q  $ (!Xd_0__inst_mult_10_27_q  $ (((Xd_0__inst_mult_10_24_q  & Xd_0__inst_mult_10_25_q )))) ) + ( Xd_0__inst_mult_10_222  ) + ( Xd_0__inst_mult_10_221  ))
// Xd_0__inst_mult_10_225  = CARRY(( !Xd_0__inst_mult_10_26_q  $ (!Xd_0__inst_mult_10_27_q  $ (((Xd_0__inst_mult_10_24_q  & Xd_0__inst_mult_10_25_q )))) ) + ( Xd_0__inst_mult_10_222  ) + ( Xd_0__inst_mult_10_221  ))
// Xd_0__inst_mult_10_226  = SHARE((Xd_0__inst_mult_10_24_q  & (Xd_0__inst_mult_10_25_q  & (!Xd_0__inst_mult_10_26_q  $ (!Xd_0__inst_mult_10_27_q )))))

	.dataa(!Xd_0__inst_mult_10_26_q ),
	.datab(!Xd_0__inst_mult_10_27_q ),
	.datac(!Xd_0__inst_mult_10_24_q ),
	.datad(!Xd_0__inst_mult_10_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_221 ),
	.sharein(Xd_0__inst_mult_10_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_224 ),
	.cout(Xd_0__inst_mult_10_225 ),
	.shareout(Xd_0__inst_mult_10_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_82 (
// Equation(s):
// Xd_0__inst_mult_11_228  = SUM(( !Xd_0__inst_mult_11_26_q  $ (!Xd_0__inst_mult_11_27_q  $ (((Xd_0__inst_mult_11_24_q  & Xd_0__inst_mult_11_25_q )))) ) + ( Xd_0__inst_mult_11_226  ) + ( Xd_0__inst_mult_11_225  ))
// Xd_0__inst_mult_11_229  = CARRY(( !Xd_0__inst_mult_11_26_q  $ (!Xd_0__inst_mult_11_27_q  $ (((Xd_0__inst_mult_11_24_q  & Xd_0__inst_mult_11_25_q )))) ) + ( Xd_0__inst_mult_11_226  ) + ( Xd_0__inst_mult_11_225  ))
// Xd_0__inst_mult_11_230  = SHARE((Xd_0__inst_mult_11_24_q  & (Xd_0__inst_mult_11_25_q  & (!Xd_0__inst_mult_11_26_q  $ (!Xd_0__inst_mult_11_27_q )))))

	.dataa(!Xd_0__inst_mult_11_26_q ),
	.datab(!Xd_0__inst_mult_11_27_q ),
	.datac(!Xd_0__inst_mult_11_24_q ),
	.datad(!Xd_0__inst_mult_11_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_225 ),
	.sharein(Xd_0__inst_mult_11_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_228 ),
	.cout(Xd_0__inst_mult_11_229 ),
	.shareout(Xd_0__inst_mult_11_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_82 (
// Equation(s):
// Xd_0__inst_mult_8_228  = SUM(( !Xd_0__inst_mult_8_26_q  $ (!Xd_0__inst_mult_8_27_q  $ (((Xd_0__inst_mult_8_24_q  & Xd_0__inst_mult_8_25_q )))) ) + ( Xd_0__inst_mult_8_226  ) + ( Xd_0__inst_mult_8_225  ))
// Xd_0__inst_mult_8_229  = CARRY(( !Xd_0__inst_mult_8_26_q  $ (!Xd_0__inst_mult_8_27_q  $ (((Xd_0__inst_mult_8_24_q  & Xd_0__inst_mult_8_25_q )))) ) + ( Xd_0__inst_mult_8_226  ) + ( Xd_0__inst_mult_8_225  ))
// Xd_0__inst_mult_8_230  = SHARE((Xd_0__inst_mult_8_24_q  & (Xd_0__inst_mult_8_25_q  & (!Xd_0__inst_mult_8_26_q  $ (!Xd_0__inst_mult_8_27_q )))))

	.dataa(!Xd_0__inst_mult_8_26_q ),
	.datab(!Xd_0__inst_mult_8_27_q ),
	.datac(!Xd_0__inst_mult_8_24_q ),
	.datad(!Xd_0__inst_mult_8_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_225 ),
	.sharein(Xd_0__inst_mult_8_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_228 ),
	.cout(Xd_0__inst_mult_8_229 ),
	.shareout(Xd_0__inst_mult_8_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_78 (
// Equation(s):
// Xd_0__inst_mult_9_224  = SUM(( !Xd_0__inst_mult_9_26_q  $ (!Xd_0__inst_mult_9_27_q  $ (((Xd_0__inst_mult_9_24_q  & Xd_0__inst_mult_9_25_q )))) ) + ( Xd_0__inst_mult_9_222  ) + ( Xd_0__inst_mult_9_221  ))
// Xd_0__inst_mult_9_225  = CARRY(( !Xd_0__inst_mult_9_26_q  $ (!Xd_0__inst_mult_9_27_q  $ (((Xd_0__inst_mult_9_24_q  & Xd_0__inst_mult_9_25_q )))) ) + ( Xd_0__inst_mult_9_222  ) + ( Xd_0__inst_mult_9_221  ))
// Xd_0__inst_mult_9_226  = SHARE((Xd_0__inst_mult_9_24_q  & (Xd_0__inst_mult_9_25_q  & (!Xd_0__inst_mult_9_26_q  $ (!Xd_0__inst_mult_9_27_q )))))

	.dataa(!Xd_0__inst_mult_9_26_q ),
	.datab(!Xd_0__inst_mult_9_27_q ),
	.datac(!Xd_0__inst_mult_9_24_q ),
	.datad(!Xd_0__inst_mult_9_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_221 ),
	.sharein(Xd_0__inst_mult_9_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_224 ),
	.cout(Xd_0__inst_mult_9_225 ),
	.shareout(Xd_0__inst_mult_9_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_78 (
// Equation(s):
// Xd_0__inst_mult_6_224  = SUM(( !Xd_0__inst_mult_6_26_q  $ (!Xd_0__inst_mult_6_27_q  $ (((Xd_0__inst_mult_6_24_q  & Xd_0__inst_mult_6_25_q )))) ) + ( Xd_0__inst_mult_6_222  ) + ( Xd_0__inst_mult_6_221  ))
// Xd_0__inst_mult_6_225  = CARRY(( !Xd_0__inst_mult_6_26_q  $ (!Xd_0__inst_mult_6_27_q  $ (((Xd_0__inst_mult_6_24_q  & Xd_0__inst_mult_6_25_q )))) ) + ( Xd_0__inst_mult_6_222  ) + ( Xd_0__inst_mult_6_221  ))
// Xd_0__inst_mult_6_226  = SHARE((Xd_0__inst_mult_6_24_q  & (Xd_0__inst_mult_6_25_q  & (!Xd_0__inst_mult_6_26_q  $ (!Xd_0__inst_mult_6_27_q )))))

	.dataa(!Xd_0__inst_mult_6_26_q ),
	.datab(!Xd_0__inst_mult_6_27_q ),
	.datac(!Xd_0__inst_mult_6_24_q ),
	.datad(!Xd_0__inst_mult_6_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_221 ),
	.sharein(Xd_0__inst_mult_6_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_224 ),
	.cout(Xd_0__inst_mult_6_225 ),
	.shareout(Xd_0__inst_mult_6_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_76 (
// Equation(s):
// Xd_0__inst_mult_7_216  = SUM(( !Xd_0__inst_mult_7_26_q  $ (!Xd_0__inst_mult_7_27_q  $ (((Xd_0__inst_mult_7_24_q  & Xd_0__inst_mult_7_25_q )))) ) + ( Xd_0__inst_mult_7_214  ) + ( Xd_0__inst_mult_7_213  ))
// Xd_0__inst_mult_7_217  = CARRY(( !Xd_0__inst_mult_7_26_q  $ (!Xd_0__inst_mult_7_27_q  $ (((Xd_0__inst_mult_7_24_q  & Xd_0__inst_mult_7_25_q )))) ) + ( Xd_0__inst_mult_7_214  ) + ( Xd_0__inst_mult_7_213  ))
// Xd_0__inst_mult_7_218  = SHARE((Xd_0__inst_mult_7_24_q  & (Xd_0__inst_mult_7_25_q  & (!Xd_0__inst_mult_7_26_q  $ (!Xd_0__inst_mult_7_27_q )))))

	.dataa(!Xd_0__inst_mult_7_26_q ),
	.datab(!Xd_0__inst_mult_7_27_q ),
	.datac(!Xd_0__inst_mult_7_24_q ),
	.datad(!Xd_0__inst_mult_7_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_213 ),
	.sharein(Xd_0__inst_mult_7_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_216 ),
	.cout(Xd_0__inst_mult_7_217 ),
	.shareout(Xd_0__inst_mult_7_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_86 (
// Equation(s):
// Xd_0__inst_mult_4_244  = SUM(( !Xd_0__inst_mult_4_26_q  $ (!Xd_0__inst_mult_4_27_q  $ (((Xd_0__inst_mult_4_24_q  & Xd_0__inst_mult_4_25_q )))) ) + ( Xd_0__inst_mult_4_242  ) + ( Xd_0__inst_mult_4_241  ))
// Xd_0__inst_mult_4_245  = CARRY(( !Xd_0__inst_mult_4_26_q  $ (!Xd_0__inst_mult_4_27_q  $ (((Xd_0__inst_mult_4_24_q  & Xd_0__inst_mult_4_25_q )))) ) + ( Xd_0__inst_mult_4_242  ) + ( Xd_0__inst_mult_4_241  ))
// Xd_0__inst_mult_4_246  = SHARE((Xd_0__inst_mult_4_24_q  & (Xd_0__inst_mult_4_25_q  & (!Xd_0__inst_mult_4_26_q  $ (!Xd_0__inst_mult_4_27_q )))))

	.dataa(!Xd_0__inst_mult_4_26_q ),
	.datab(!Xd_0__inst_mult_4_27_q ),
	.datac(!Xd_0__inst_mult_4_24_q ),
	.datad(!Xd_0__inst_mult_4_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_241 ),
	.sharein(Xd_0__inst_mult_4_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_244 ),
	.cout(Xd_0__inst_mult_4_245 ),
	.shareout(Xd_0__inst_mult_4_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_76 (
// Equation(s):
// Xd_0__inst_mult_5_216  = SUM(( !Xd_0__inst_mult_5_26_q  $ (!Xd_0__inst_mult_5_27_q  $ (((Xd_0__inst_mult_5_24_q  & Xd_0__inst_mult_5_25_q )))) ) + ( Xd_0__inst_mult_5_214  ) + ( Xd_0__inst_mult_5_213  ))
// Xd_0__inst_mult_5_217  = CARRY(( !Xd_0__inst_mult_5_26_q  $ (!Xd_0__inst_mult_5_27_q  $ (((Xd_0__inst_mult_5_24_q  & Xd_0__inst_mult_5_25_q )))) ) + ( Xd_0__inst_mult_5_214  ) + ( Xd_0__inst_mult_5_213  ))
// Xd_0__inst_mult_5_218  = SHARE((Xd_0__inst_mult_5_24_q  & (Xd_0__inst_mult_5_25_q  & (!Xd_0__inst_mult_5_26_q  $ (!Xd_0__inst_mult_5_27_q )))))

	.dataa(!Xd_0__inst_mult_5_26_q ),
	.datab(!Xd_0__inst_mult_5_27_q ),
	.datac(!Xd_0__inst_mult_5_24_q ),
	.datad(!Xd_0__inst_mult_5_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_213 ),
	.sharein(Xd_0__inst_mult_5_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_216 ),
	.cout(Xd_0__inst_mult_5_217 ),
	.shareout(Xd_0__inst_mult_5_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_80 (
// Equation(s):
// Xd_0__inst_mult_2_220  = SUM(( !Xd_0__inst_mult_2_26_q  $ (!Xd_0__inst_mult_2_27_q  $ (((Xd_0__inst_mult_2_24_q  & Xd_0__inst_mult_2_25_q )))) ) + ( Xd_0__inst_mult_2_218  ) + ( Xd_0__inst_mult_2_217  ))
// Xd_0__inst_mult_2_221  = CARRY(( !Xd_0__inst_mult_2_26_q  $ (!Xd_0__inst_mult_2_27_q  $ (((Xd_0__inst_mult_2_24_q  & Xd_0__inst_mult_2_25_q )))) ) + ( Xd_0__inst_mult_2_218  ) + ( Xd_0__inst_mult_2_217  ))
// Xd_0__inst_mult_2_222  = SHARE((Xd_0__inst_mult_2_24_q  & (Xd_0__inst_mult_2_25_q  & (!Xd_0__inst_mult_2_26_q  $ (!Xd_0__inst_mult_2_27_q )))))

	.dataa(!Xd_0__inst_mult_2_26_q ),
	.datab(!Xd_0__inst_mult_2_27_q ),
	.datac(!Xd_0__inst_mult_2_24_q ),
	.datad(!Xd_0__inst_mult_2_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_217 ),
	.sharein(Xd_0__inst_mult_2_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_220 ),
	.cout(Xd_0__inst_mult_2_221 ),
	.shareout(Xd_0__inst_mult_2_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_76 (
// Equation(s):
// Xd_0__inst_mult_3_216  = SUM(( !Xd_0__inst_mult_3_26_q  $ (!Xd_0__inst_mult_3_27_q  $ (((Xd_0__inst_mult_3_24_q  & Xd_0__inst_mult_3_25_q )))) ) + ( Xd_0__inst_mult_3_214  ) + ( Xd_0__inst_mult_3_213  ))
// Xd_0__inst_mult_3_217  = CARRY(( !Xd_0__inst_mult_3_26_q  $ (!Xd_0__inst_mult_3_27_q  $ (((Xd_0__inst_mult_3_24_q  & Xd_0__inst_mult_3_25_q )))) ) + ( Xd_0__inst_mult_3_214  ) + ( Xd_0__inst_mult_3_213  ))
// Xd_0__inst_mult_3_218  = SHARE((Xd_0__inst_mult_3_24_q  & (Xd_0__inst_mult_3_25_q  & (!Xd_0__inst_mult_3_26_q  $ (!Xd_0__inst_mult_3_27_q )))))

	.dataa(!Xd_0__inst_mult_3_26_q ),
	.datab(!Xd_0__inst_mult_3_27_q ),
	.datac(!Xd_0__inst_mult_3_24_q ),
	.datad(!Xd_0__inst_mult_3_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_213 ),
	.sharein(Xd_0__inst_mult_3_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_216 ),
	.cout(Xd_0__inst_mult_3_217 ),
	.shareout(Xd_0__inst_mult_3_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_80 (
// Equation(s):
// Xd_0__inst_mult_0_220  = SUM(( !Xd_0__inst_mult_0_26_q  $ (!Xd_0__inst_mult_0_27_q  $ (((Xd_0__inst_mult_0_24_q  & Xd_0__inst_mult_0_25_q )))) ) + ( Xd_0__inst_mult_0_218  ) + ( Xd_0__inst_mult_0_217  ))
// Xd_0__inst_mult_0_221  = CARRY(( !Xd_0__inst_mult_0_26_q  $ (!Xd_0__inst_mult_0_27_q  $ (((Xd_0__inst_mult_0_24_q  & Xd_0__inst_mult_0_25_q )))) ) + ( Xd_0__inst_mult_0_218  ) + ( Xd_0__inst_mult_0_217  ))
// Xd_0__inst_mult_0_222  = SHARE((Xd_0__inst_mult_0_24_q  & (Xd_0__inst_mult_0_25_q  & (!Xd_0__inst_mult_0_26_q  $ (!Xd_0__inst_mult_0_27_q )))))

	.dataa(!Xd_0__inst_mult_0_26_q ),
	.datab(!Xd_0__inst_mult_0_27_q ),
	.datac(!Xd_0__inst_mult_0_24_q ),
	.datad(!Xd_0__inst_mult_0_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_217 ),
	.sharein(Xd_0__inst_mult_0_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_220 ),
	.cout(Xd_0__inst_mult_0_221 ),
	.shareout(Xd_0__inst_mult_0_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_80 (
// Equation(s):
// Xd_0__inst_mult_1_220  = SUM(( !Xd_0__inst_mult_1_26_q  $ (!Xd_0__inst_mult_1_27_q  $ (((Xd_0__inst_mult_1_24_q  & Xd_0__inst_mult_1_25_q )))) ) + ( Xd_0__inst_mult_1_218  ) + ( Xd_0__inst_mult_1_217  ))
// Xd_0__inst_mult_1_221  = CARRY(( !Xd_0__inst_mult_1_26_q  $ (!Xd_0__inst_mult_1_27_q  $ (((Xd_0__inst_mult_1_24_q  & Xd_0__inst_mult_1_25_q )))) ) + ( Xd_0__inst_mult_1_218  ) + ( Xd_0__inst_mult_1_217  ))
// Xd_0__inst_mult_1_222  = SHARE((Xd_0__inst_mult_1_24_q  & (Xd_0__inst_mult_1_25_q  & (!Xd_0__inst_mult_1_26_q  $ (!Xd_0__inst_mult_1_27_q )))))

	.dataa(!Xd_0__inst_mult_1_26_q ),
	.datab(!Xd_0__inst_mult_1_27_q ),
	.datac(!Xd_0__inst_mult_1_24_q ),
	.datad(!Xd_0__inst_mult_1_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_217 ),
	.sharein(Xd_0__inst_mult_1_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_220 ),
	.cout(Xd_0__inst_mult_1_221 ),
	.shareout(Xd_0__inst_mult_1_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_83 (
// Equation(s):
// Xd_0__inst_mult_12_244  = SUM(( !Xd_0__inst_mult_12_28_q  $ (!Xd_0__inst_mult_12_29_q  $ (((Xd_0__inst_mult_12_26_q  & Xd_0__inst_mult_12_27_q )))) ) + ( Xd_0__inst_mult_12_242  ) + ( Xd_0__inst_mult_12_241  ))
// Xd_0__inst_mult_12_245  = CARRY(( !Xd_0__inst_mult_12_28_q  $ (!Xd_0__inst_mult_12_29_q  $ (((Xd_0__inst_mult_12_26_q  & Xd_0__inst_mult_12_27_q )))) ) + ( Xd_0__inst_mult_12_242  ) + ( Xd_0__inst_mult_12_241  ))
// Xd_0__inst_mult_12_246  = SHARE((Xd_0__inst_mult_12_26_q  & (Xd_0__inst_mult_12_27_q  & (!Xd_0__inst_mult_12_28_q  $ (!Xd_0__inst_mult_12_29_q )))))

	.dataa(!Xd_0__inst_mult_12_28_q ),
	.datab(!Xd_0__inst_mult_12_29_q ),
	.datac(!Xd_0__inst_mult_12_26_q ),
	.datad(!Xd_0__inst_mult_12_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_241 ),
	.sharein(Xd_0__inst_mult_12_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_244 ),
	.cout(Xd_0__inst_mult_12_245 ),
	.shareout(Xd_0__inst_mult_12_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_83 (
// Equation(s):
// Xd_0__inst_mult_13_232  = SUM(( !Xd_0__inst_mult_13_28_q  $ (!Xd_0__inst_mult_13_29_q  $ (((Xd_0__inst_mult_13_26_q  & Xd_0__inst_mult_13_27_q )))) ) + ( Xd_0__inst_mult_13_230  ) + ( Xd_0__inst_mult_13_229  ))
// Xd_0__inst_mult_13_233  = CARRY(( !Xd_0__inst_mult_13_28_q  $ (!Xd_0__inst_mult_13_29_q  $ (((Xd_0__inst_mult_13_26_q  & Xd_0__inst_mult_13_27_q )))) ) + ( Xd_0__inst_mult_13_230  ) + ( Xd_0__inst_mult_13_229  ))
// Xd_0__inst_mult_13_234  = SHARE((Xd_0__inst_mult_13_26_q  & (Xd_0__inst_mult_13_27_q  & (!Xd_0__inst_mult_13_28_q  $ (!Xd_0__inst_mult_13_29_q )))))

	.dataa(!Xd_0__inst_mult_13_28_q ),
	.datab(!Xd_0__inst_mult_13_29_q ),
	.datac(!Xd_0__inst_mult_13_26_q ),
	.datad(!Xd_0__inst_mult_13_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_229 ),
	.sharein(Xd_0__inst_mult_13_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_232 ),
	.cout(Xd_0__inst_mult_13_233 ),
	.shareout(Xd_0__inst_mult_13_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_87 (
// Equation(s):
// Xd_0__inst_mult_14_248  = SUM(( !Xd_0__inst_mult_14_28_q  $ (!Xd_0__inst_mult_14_29_q  $ (((Xd_0__inst_mult_14_26_q  & Xd_0__inst_mult_14_27_q )))) ) + ( Xd_0__inst_mult_14_246  ) + ( Xd_0__inst_mult_14_245  ))
// Xd_0__inst_mult_14_249  = CARRY(( !Xd_0__inst_mult_14_28_q  $ (!Xd_0__inst_mult_14_29_q  $ (((Xd_0__inst_mult_14_26_q  & Xd_0__inst_mult_14_27_q )))) ) + ( Xd_0__inst_mult_14_246  ) + ( Xd_0__inst_mult_14_245  ))
// Xd_0__inst_mult_14_250  = SHARE((Xd_0__inst_mult_14_26_q  & (Xd_0__inst_mult_14_27_q  & (!Xd_0__inst_mult_14_28_q  $ (!Xd_0__inst_mult_14_29_q )))))

	.dataa(!Xd_0__inst_mult_14_28_q ),
	.datab(!Xd_0__inst_mult_14_29_q ),
	.datac(!Xd_0__inst_mult_14_26_q ),
	.datad(!Xd_0__inst_mult_14_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_245 ),
	.sharein(Xd_0__inst_mult_14_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_248 ),
	.cout(Xd_0__inst_mult_14_249 ),
	.shareout(Xd_0__inst_mult_14_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_87 (
// Equation(s):
// Xd_0__inst_mult_15_248  = SUM(( !Xd_0__inst_mult_15_28_q  $ (!Xd_0__inst_mult_15_29_q  $ (((Xd_0__inst_mult_15_26_q  & Xd_0__inst_mult_15_27_q )))) ) + ( Xd_0__inst_mult_15_246  ) + ( Xd_0__inst_mult_15_245  ))
// Xd_0__inst_mult_15_249  = CARRY(( !Xd_0__inst_mult_15_28_q  $ (!Xd_0__inst_mult_15_29_q  $ (((Xd_0__inst_mult_15_26_q  & Xd_0__inst_mult_15_27_q )))) ) + ( Xd_0__inst_mult_15_246  ) + ( Xd_0__inst_mult_15_245  ))
// Xd_0__inst_mult_15_250  = SHARE((Xd_0__inst_mult_15_26_q  & (Xd_0__inst_mult_15_27_q  & (!Xd_0__inst_mult_15_28_q  $ (!Xd_0__inst_mult_15_29_q )))))

	.dataa(!Xd_0__inst_mult_15_28_q ),
	.datab(!Xd_0__inst_mult_15_29_q ),
	.datac(!Xd_0__inst_mult_15_26_q ),
	.datad(!Xd_0__inst_mult_15_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_245 ),
	.sharein(Xd_0__inst_mult_15_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_248 ),
	.cout(Xd_0__inst_mult_15_249 ),
	.shareout(Xd_0__inst_mult_15_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_79 (
// Equation(s):
// Xd_0__inst_mult_10_228  = SUM(( !Xd_0__inst_mult_10_28_q  $ (!Xd_0__inst_mult_10_29_q  $ (((Xd_0__inst_mult_10_26_q  & Xd_0__inst_mult_10_27_q )))) ) + ( Xd_0__inst_mult_10_226  ) + ( Xd_0__inst_mult_10_225  ))
// Xd_0__inst_mult_10_229  = CARRY(( !Xd_0__inst_mult_10_28_q  $ (!Xd_0__inst_mult_10_29_q  $ (((Xd_0__inst_mult_10_26_q  & Xd_0__inst_mult_10_27_q )))) ) + ( Xd_0__inst_mult_10_226  ) + ( Xd_0__inst_mult_10_225  ))
// Xd_0__inst_mult_10_230  = SHARE((Xd_0__inst_mult_10_26_q  & (Xd_0__inst_mult_10_27_q  & (!Xd_0__inst_mult_10_28_q  $ (!Xd_0__inst_mult_10_29_q )))))

	.dataa(!Xd_0__inst_mult_10_28_q ),
	.datab(!Xd_0__inst_mult_10_29_q ),
	.datac(!Xd_0__inst_mult_10_26_q ),
	.datad(!Xd_0__inst_mult_10_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_225 ),
	.sharein(Xd_0__inst_mult_10_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_228 ),
	.cout(Xd_0__inst_mult_10_229 ),
	.shareout(Xd_0__inst_mult_10_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_83 (
// Equation(s):
// Xd_0__inst_mult_11_232  = SUM(( !Xd_0__inst_mult_11_28_q  $ (!Xd_0__inst_mult_11_29_q  $ (((Xd_0__inst_mult_11_26_q  & Xd_0__inst_mult_11_27_q )))) ) + ( Xd_0__inst_mult_11_230  ) + ( Xd_0__inst_mult_11_229  ))
// Xd_0__inst_mult_11_233  = CARRY(( !Xd_0__inst_mult_11_28_q  $ (!Xd_0__inst_mult_11_29_q  $ (((Xd_0__inst_mult_11_26_q  & Xd_0__inst_mult_11_27_q )))) ) + ( Xd_0__inst_mult_11_230  ) + ( Xd_0__inst_mult_11_229  ))
// Xd_0__inst_mult_11_234  = SHARE((Xd_0__inst_mult_11_26_q  & (Xd_0__inst_mult_11_27_q  & (!Xd_0__inst_mult_11_28_q  $ (!Xd_0__inst_mult_11_29_q )))))

	.dataa(!Xd_0__inst_mult_11_28_q ),
	.datab(!Xd_0__inst_mult_11_29_q ),
	.datac(!Xd_0__inst_mult_11_26_q ),
	.datad(!Xd_0__inst_mult_11_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_229 ),
	.sharein(Xd_0__inst_mult_11_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_232 ),
	.cout(Xd_0__inst_mult_11_233 ),
	.shareout(Xd_0__inst_mult_11_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_83 (
// Equation(s):
// Xd_0__inst_mult_8_232  = SUM(( !Xd_0__inst_mult_8_28_q  $ (!Xd_0__inst_mult_8_29_q  $ (((Xd_0__inst_mult_8_26_q  & Xd_0__inst_mult_8_27_q )))) ) + ( Xd_0__inst_mult_8_230  ) + ( Xd_0__inst_mult_8_229  ))
// Xd_0__inst_mult_8_233  = CARRY(( !Xd_0__inst_mult_8_28_q  $ (!Xd_0__inst_mult_8_29_q  $ (((Xd_0__inst_mult_8_26_q  & Xd_0__inst_mult_8_27_q )))) ) + ( Xd_0__inst_mult_8_230  ) + ( Xd_0__inst_mult_8_229  ))
// Xd_0__inst_mult_8_234  = SHARE((Xd_0__inst_mult_8_26_q  & (Xd_0__inst_mult_8_27_q  & (!Xd_0__inst_mult_8_28_q  $ (!Xd_0__inst_mult_8_29_q )))))

	.dataa(!Xd_0__inst_mult_8_28_q ),
	.datab(!Xd_0__inst_mult_8_29_q ),
	.datac(!Xd_0__inst_mult_8_26_q ),
	.datad(!Xd_0__inst_mult_8_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_229 ),
	.sharein(Xd_0__inst_mult_8_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_232 ),
	.cout(Xd_0__inst_mult_8_233 ),
	.shareout(Xd_0__inst_mult_8_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_79 (
// Equation(s):
// Xd_0__inst_mult_9_228  = SUM(( !Xd_0__inst_mult_9_28_q  $ (!Xd_0__inst_mult_9_29_q  $ (((Xd_0__inst_mult_9_26_q  & Xd_0__inst_mult_9_27_q )))) ) + ( Xd_0__inst_mult_9_226  ) + ( Xd_0__inst_mult_9_225  ))
// Xd_0__inst_mult_9_229  = CARRY(( !Xd_0__inst_mult_9_28_q  $ (!Xd_0__inst_mult_9_29_q  $ (((Xd_0__inst_mult_9_26_q  & Xd_0__inst_mult_9_27_q )))) ) + ( Xd_0__inst_mult_9_226  ) + ( Xd_0__inst_mult_9_225  ))
// Xd_0__inst_mult_9_230  = SHARE((Xd_0__inst_mult_9_26_q  & (Xd_0__inst_mult_9_27_q  & (!Xd_0__inst_mult_9_28_q  $ (!Xd_0__inst_mult_9_29_q )))))

	.dataa(!Xd_0__inst_mult_9_28_q ),
	.datab(!Xd_0__inst_mult_9_29_q ),
	.datac(!Xd_0__inst_mult_9_26_q ),
	.datad(!Xd_0__inst_mult_9_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_225 ),
	.sharein(Xd_0__inst_mult_9_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_228 ),
	.cout(Xd_0__inst_mult_9_229 ),
	.shareout(Xd_0__inst_mult_9_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_79 (
// Equation(s):
// Xd_0__inst_mult_6_228  = SUM(( !Xd_0__inst_mult_6_28_q  $ (!Xd_0__inst_mult_6_29_q  $ (((Xd_0__inst_mult_6_26_q  & Xd_0__inst_mult_6_27_q )))) ) + ( Xd_0__inst_mult_6_226  ) + ( Xd_0__inst_mult_6_225  ))
// Xd_0__inst_mult_6_229  = CARRY(( !Xd_0__inst_mult_6_28_q  $ (!Xd_0__inst_mult_6_29_q  $ (((Xd_0__inst_mult_6_26_q  & Xd_0__inst_mult_6_27_q )))) ) + ( Xd_0__inst_mult_6_226  ) + ( Xd_0__inst_mult_6_225  ))
// Xd_0__inst_mult_6_230  = SHARE((Xd_0__inst_mult_6_26_q  & (Xd_0__inst_mult_6_27_q  & (!Xd_0__inst_mult_6_28_q  $ (!Xd_0__inst_mult_6_29_q )))))

	.dataa(!Xd_0__inst_mult_6_28_q ),
	.datab(!Xd_0__inst_mult_6_29_q ),
	.datac(!Xd_0__inst_mult_6_26_q ),
	.datad(!Xd_0__inst_mult_6_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_225 ),
	.sharein(Xd_0__inst_mult_6_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_228 ),
	.cout(Xd_0__inst_mult_6_229 ),
	.shareout(Xd_0__inst_mult_6_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_77 (
// Equation(s):
// Xd_0__inst_mult_7_220  = SUM(( !Xd_0__inst_mult_7_28_q  $ (!Xd_0__inst_mult_7_29_q  $ (((Xd_0__inst_mult_7_26_q  & Xd_0__inst_mult_7_27_q )))) ) + ( Xd_0__inst_mult_7_218  ) + ( Xd_0__inst_mult_7_217  ))
// Xd_0__inst_mult_7_221  = CARRY(( !Xd_0__inst_mult_7_28_q  $ (!Xd_0__inst_mult_7_29_q  $ (((Xd_0__inst_mult_7_26_q  & Xd_0__inst_mult_7_27_q )))) ) + ( Xd_0__inst_mult_7_218  ) + ( Xd_0__inst_mult_7_217  ))
// Xd_0__inst_mult_7_222  = SHARE((Xd_0__inst_mult_7_26_q  & (Xd_0__inst_mult_7_27_q  & (!Xd_0__inst_mult_7_28_q  $ (!Xd_0__inst_mult_7_29_q )))))

	.dataa(!Xd_0__inst_mult_7_28_q ),
	.datab(!Xd_0__inst_mult_7_29_q ),
	.datac(!Xd_0__inst_mult_7_26_q ),
	.datad(!Xd_0__inst_mult_7_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_217 ),
	.sharein(Xd_0__inst_mult_7_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_220 ),
	.cout(Xd_0__inst_mult_7_221 ),
	.shareout(Xd_0__inst_mult_7_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_87 (
// Equation(s):
// Xd_0__inst_mult_4_248  = SUM(( !Xd_0__inst_mult_4_28_q  $ (!Xd_0__inst_mult_4_29_q  $ (((Xd_0__inst_mult_4_26_q  & Xd_0__inst_mult_4_27_q )))) ) + ( Xd_0__inst_mult_4_246  ) + ( Xd_0__inst_mult_4_245  ))
// Xd_0__inst_mult_4_249  = CARRY(( !Xd_0__inst_mult_4_28_q  $ (!Xd_0__inst_mult_4_29_q  $ (((Xd_0__inst_mult_4_26_q  & Xd_0__inst_mult_4_27_q )))) ) + ( Xd_0__inst_mult_4_246  ) + ( Xd_0__inst_mult_4_245  ))
// Xd_0__inst_mult_4_250  = SHARE((Xd_0__inst_mult_4_26_q  & (Xd_0__inst_mult_4_27_q  & (!Xd_0__inst_mult_4_28_q  $ (!Xd_0__inst_mult_4_29_q )))))

	.dataa(!Xd_0__inst_mult_4_28_q ),
	.datab(!Xd_0__inst_mult_4_29_q ),
	.datac(!Xd_0__inst_mult_4_26_q ),
	.datad(!Xd_0__inst_mult_4_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_245 ),
	.sharein(Xd_0__inst_mult_4_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_248 ),
	.cout(Xd_0__inst_mult_4_249 ),
	.shareout(Xd_0__inst_mult_4_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_77 (
// Equation(s):
// Xd_0__inst_mult_5_220  = SUM(( !Xd_0__inst_mult_5_28_q  $ (!Xd_0__inst_mult_5_29_q  $ (((Xd_0__inst_mult_5_26_q  & Xd_0__inst_mult_5_27_q )))) ) + ( Xd_0__inst_mult_5_218  ) + ( Xd_0__inst_mult_5_217  ))
// Xd_0__inst_mult_5_221  = CARRY(( !Xd_0__inst_mult_5_28_q  $ (!Xd_0__inst_mult_5_29_q  $ (((Xd_0__inst_mult_5_26_q  & Xd_0__inst_mult_5_27_q )))) ) + ( Xd_0__inst_mult_5_218  ) + ( Xd_0__inst_mult_5_217  ))
// Xd_0__inst_mult_5_222  = SHARE((Xd_0__inst_mult_5_26_q  & (Xd_0__inst_mult_5_27_q  & (!Xd_0__inst_mult_5_28_q  $ (!Xd_0__inst_mult_5_29_q )))))

	.dataa(!Xd_0__inst_mult_5_28_q ),
	.datab(!Xd_0__inst_mult_5_29_q ),
	.datac(!Xd_0__inst_mult_5_26_q ),
	.datad(!Xd_0__inst_mult_5_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_217 ),
	.sharein(Xd_0__inst_mult_5_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_220 ),
	.cout(Xd_0__inst_mult_5_221 ),
	.shareout(Xd_0__inst_mult_5_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_81 (
// Equation(s):
// Xd_0__inst_mult_2_224  = SUM(( !Xd_0__inst_mult_2_28_q  $ (!Xd_0__inst_mult_2_29_q  $ (((Xd_0__inst_mult_2_26_q  & Xd_0__inst_mult_2_27_q )))) ) + ( Xd_0__inst_mult_2_222  ) + ( Xd_0__inst_mult_2_221  ))
// Xd_0__inst_mult_2_225  = CARRY(( !Xd_0__inst_mult_2_28_q  $ (!Xd_0__inst_mult_2_29_q  $ (((Xd_0__inst_mult_2_26_q  & Xd_0__inst_mult_2_27_q )))) ) + ( Xd_0__inst_mult_2_222  ) + ( Xd_0__inst_mult_2_221  ))
// Xd_0__inst_mult_2_226  = SHARE((Xd_0__inst_mult_2_26_q  & (Xd_0__inst_mult_2_27_q  & (!Xd_0__inst_mult_2_28_q  $ (!Xd_0__inst_mult_2_29_q )))))

	.dataa(!Xd_0__inst_mult_2_28_q ),
	.datab(!Xd_0__inst_mult_2_29_q ),
	.datac(!Xd_0__inst_mult_2_26_q ),
	.datad(!Xd_0__inst_mult_2_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_221 ),
	.sharein(Xd_0__inst_mult_2_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_224 ),
	.cout(Xd_0__inst_mult_2_225 ),
	.shareout(Xd_0__inst_mult_2_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_77 (
// Equation(s):
// Xd_0__inst_mult_3_220  = SUM(( !Xd_0__inst_mult_3_28_q  $ (!Xd_0__inst_mult_3_29_q  $ (((Xd_0__inst_mult_3_26_q  & Xd_0__inst_mult_3_27_q )))) ) + ( Xd_0__inst_mult_3_218  ) + ( Xd_0__inst_mult_3_217  ))
// Xd_0__inst_mult_3_221  = CARRY(( !Xd_0__inst_mult_3_28_q  $ (!Xd_0__inst_mult_3_29_q  $ (((Xd_0__inst_mult_3_26_q  & Xd_0__inst_mult_3_27_q )))) ) + ( Xd_0__inst_mult_3_218  ) + ( Xd_0__inst_mult_3_217  ))
// Xd_0__inst_mult_3_222  = SHARE((Xd_0__inst_mult_3_26_q  & (Xd_0__inst_mult_3_27_q  & (!Xd_0__inst_mult_3_28_q  $ (!Xd_0__inst_mult_3_29_q )))))

	.dataa(!Xd_0__inst_mult_3_28_q ),
	.datab(!Xd_0__inst_mult_3_29_q ),
	.datac(!Xd_0__inst_mult_3_26_q ),
	.datad(!Xd_0__inst_mult_3_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_217 ),
	.sharein(Xd_0__inst_mult_3_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_220 ),
	.cout(Xd_0__inst_mult_3_221 ),
	.shareout(Xd_0__inst_mult_3_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_81 (
// Equation(s):
// Xd_0__inst_mult_0_224  = SUM(( !Xd_0__inst_mult_0_28_q  $ (!Xd_0__inst_mult_0_29_q  $ (((Xd_0__inst_mult_0_26_q  & Xd_0__inst_mult_0_27_q )))) ) + ( Xd_0__inst_mult_0_222  ) + ( Xd_0__inst_mult_0_221  ))
// Xd_0__inst_mult_0_225  = CARRY(( !Xd_0__inst_mult_0_28_q  $ (!Xd_0__inst_mult_0_29_q  $ (((Xd_0__inst_mult_0_26_q  & Xd_0__inst_mult_0_27_q )))) ) + ( Xd_0__inst_mult_0_222  ) + ( Xd_0__inst_mult_0_221  ))
// Xd_0__inst_mult_0_226  = SHARE((Xd_0__inst_mult_0_26_q  & (Xd_0__inst_mult_0_27_q  & (!Xd_0__inst_mult_0_28_q  $ (!Xd_0__inst_mult_0_29_q )))))

	.dataa(!Xd_0__inst_mult_0_28_q ),
	.datab(!Xd_0__inst_mult_0_29_q ),
	.datac(!Xd_0__inst_mult_0_26_q ),
	.datad(!Xd_0__inst_mult_0_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_221 ),
	.sharein(Xd_0__inst_mult_0_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_224 ),
	.cout(Xd_0__inst_mult_0_225 ),
	.shareout(Xd_0__inst_mult_0_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_81 (
// Equation(s):
// Xd_0__inst_mult_1_224  = SUM(( !Xd_0__inst_mult_1_28_q  $ (!Xd_0__inst_mult_1_29_q  $ (((Xd_0__inst_mult_1_26_q  & Xd_0__inst_mult_1_27_q )))) ) + ( Xd_0__inst_mult_1_222  ) + ( Xd_0__inst_mult_1_221  ))
// Xd_0__inst_mult_1_225  = CARRY(( !Xd_0__inst_mult_1_28_q  $ (!Xd_0__inst_mult_1_29_q  $ (((Xd_0__inst_mult_1_26_q  & Xd_0__inst_mult_1_27_q )))) ) + ( Xd_0__inst_mult_1_222  ) + ( Xd_0__inst_mult_1_221  ))
// Xd_0__inst_mult_1_226  = SHARE((Xd_0__inst_mult_1_26_q  & (Xd_0__inst_mult_1_27_q  & (!Xd_0__inst_mult_1_28_q  $ (!Xd_0__inst_mult_1_29_q )))))

	.dataa(!Xd_0__inst_mult_1_28_q ),
	.datab(!Xd_0__inst_mult_1_29_q ),
	.datac(!Xd_0__inst_mult_1_26_q ),
	.datad(!Xd_0__inst_mult_1_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_221 ),
	.sharein(Xd_0__inst_mult_1_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_224 ),
	.cout(Xd_0__inst_mult_1_225 ),
	.shareout(Xd_0__inst_mult_1_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_84 (
// Equation(s):
// Xd_0__inst_mult_12_248  = SUM(( !Xd_0__inst_mult_12_30_q  $ (!Xd_0__inst_mult_12_31_q  $ (((Xd_0__inst_mult_12_28_q  & Xd_0__inst_mult_12_29_q )))) ) + ( Xd_0__inst_mult_12_246  ) + ( Xd_0__inst_mult_12_245  ))
// Xd_0__inst_mult_12_249  = CARRY(( !Xd_0__inst_mult_12_30_q  $ (!Xd_0__inst_mult_12_31_q  $ (((Xd_0__inst_mult_12_28_q  & Xd_0__inst_mult_12_29_q )))) ) + ( Xd_0__inst_mult_12_246  ) + ( Xd_0__inst_mult_12_245  ))
// Xd_0__inst_mult_12_250  = SHARE((Xd_0__inst_mult_12_28_q  & (Xd_0__inst_mult_12_29_q  & (!Xd_0__inst_mult_12_30_q  $ (!Xd_0__inst_mult_12_31_q )))))

	.dataa(!Xd_0__inst_mult_12_30_q ),
	.datab(!Xd_0__inst_mult_12_31_q ),
	.datac(!Xd_0__inst_mult_12_28_q ),
	.datad(!Xd_0__inst_mult_12_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_245 ),
	.sharein(Xd_0__inst_mult_12_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_248 ),
	.cout(Xd_0__inst_mult_12_249 ),
	.shareout(Xd_0__inst_mult_12_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_84 (
// Equation(s):
// Xd_0__inst_mult_13_236  = SUM(( !Xd_0__inst_mult_13_30_q  $ (!Xd_0__inst_mult_13_31_q  $ (((Xd_0__inst_mult_13_28_q  & Xd_0__inst_mult_13_29_q )))) ) + ( Xd_0__inst_mult_13_234  ) + ( Xd_0__inst_mult_13_233  ))
// Xd_0__inst_mult_13_237  = CARRY(( !Xd_0__inst_mult_13_30_q  $ (!Xd_0__inst_mult_13_31_q  $ (((Xd_0__inst_mult_13_28_q  & Xd_0__inst_mult_13_29_q )))) ) + ( Xd_0__inst_mult_13_234  ) + ( Xd_0__inst_mult_13_233  ))
// Xd_0__inst_mult_13_238  = SHARE((Xd_0__inst_mult_13_28_q  & (Xd_0__inst_mult_13_29_q  & (!Xd_0__inst_mult_13_30_q  $ (!Xd_0__inst_mult_13_31_q )))))

	.dataa(!Xd_0__inst_mult_13_30_q ),
	.datab(!Xd_0__inst_mult_13_31_q ),
	.datac(!Xd_0__inst_mult_13_28_q ),
	.datad(!Xd_0__inst_mult_13_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_233 ),
	.sharein(Xd_0__inst_mult_13_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_236 ),
	.cout(Xd_0__inst_mult_13_237 ),
	.shareout(Xd_0__inst_mult_13_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_88 (
// Equation(s):
// Xd_0__inst_mult_14_252  = SUM(( !Xd_0__inst_mult_14_30_q  $ (!Xd_0__inst_mult_14_31_q  $ (((Xd_0__inst_mult_14_28_q  & Xd_0__inst_mult_14_29_q )))) ) + ( Xd_0__inst_mult_14_250  ) + ( Xd_0__inst_mult_14_249  ))
// Xd_0__inst_mult_14_253  = CARRY(( !Xd_0__inst_mult_14_30_q  $ (!Xd_0__inst_mult_14_31_q  $ (((Xd_0__inst_mult_14_28_q  & Xd_0__inst_mult_14_29_q )))) ) + ( Xd_0__inst_mult_14_250  ) + ( Xd_0__inst_mult_14_249  ))
// Xd_0__inst_mult_14_254  = SHARE((Xd_0__inst_mult_14_28_q  & (Xd_0__inst_mult_14_29_q  & (!Xd_0__inst_mult_14_30_q  $ (!Xd_0__inst_mult_14_31_q )))))

	.dataa(!Xd_0__inst_mult_14_30_q ),
	.datab(!Xd_0__inst_mult_14_31_q ),
	.datac(!Xd_0__inst_mult_14_28_q ),
	.datad(!Xd_0__inst_mult_14_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_249 ),
	.sharein(Xd_0__inst_mult_14_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_252 ),
	.cout(Xd_0__inst_mult_14_253 ),
	.shareout(Xd_0__inst_mult_14_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_88 (
// Equation(s):
// Xd_0__inst_mult_15_252  = SUM(( !Xd_0__inst_mult_15_30_q  $ (!Xd_0__inst_mult_15_31_q  $ (((Xd_0__inst_mult_15_28_q  & Xd_0__inst_mult_15_29_q )))) ) + ( Xd_0__inst_mult_15_250  ) + ( Xd_0__inst_mult_15_249  ))
// Xd_0__inst_mult_15_253  = CARRY(( !Xd_0__inst_mult_15_30_q  $ (!Xd_0__inst_mult_15_31_q  $ (((Xd_0__inst_mult_15_28_q  & Xd_0__inst_mult_15_29_q )))) ) + ( Xd_0__inst_mult_15_250  ) + ( Xd_0__inst_mult_15_249  ))
// Xd_0__inst_mult_15_254  = SHARE((Xd_0__inst_mult_15_28_q  & (Xd_0__inst_mult_15_29_q  & (!Xd_0__inst_mult_15_30_q  $ (!Xd_0__inst_mult_15_31_q )))))

	.dataa(!Xd_0__inst_mult_15_30_q ),
	.datab(!Xd_0__inst_mult_15_31_q ),
	.datac(!Xd_0__inst_mult_15_28_q ),
	.datad(!Xd_0__inst_mult_15_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_249 ),
	.sharein(Xd_0__inst_mult_15_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_252 ),
	.cout(Xd_0__inst_mult_15_253 ),
	.shareout(Xd_0__inst_mult_15_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_80 (
// Equation(s):
// Xd_0__inst_mult_10_232  = SUM(( !Xd_0__inst_mult_10_30_q  $ (!Xd_0__inst_mult_10_31_q  $ (((Xd_0__inst_mult_10_28_q  & Xd_0__inst_mult_10_29_q )))) ) + ( Xd_0__inst_mult_10_230  ) + ( Xd_0__inst_mult_10_229  ))
// Xd_0__inst_mult_10_233  = CARRY(( !Xd_0__inst_mult_10_30_q  $ (!Xd_0__inst_mult_10_31_q  $ (((Xd_0__inst_mult_10_28_q  & Xd_0__inst_mult_10_29_q )))) ) + ( Xd_0__inst_mult_10_230  ) + ( Xd_0__inst_mult_10_229  ))
// Xd_0__inst_mult_10_234  = SHARE((Xd_0__inst_mult_10_28_q  & (Xd_0__inst_mult_10_29_q  & (!Xd_0__inst_mult_10_30_q  $ (!Xd_0__inst_mult_10_31_q )))))

	.dataa(!Xd_0__inst_mult_10_30_q ),
	.datab(!Xd_0__inst_mult_10_31_q ),
	.datac(!Xd_0__inst_mult_10_28_q ),
	.datad(!Xd_0__inst_mult_10_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_229 ),
	.sharein(Xd_0__inst_mult_10_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_232 ),
	.cout(Xd_0__inst_mult_10_233 ),
	.shareout(Xd_0__inst_mult_10_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_84 (
// Equation(s):
// Xd_0__inst_mult_11_236  = SUM(( !Xd_0__inst_mult_11_30_q  $ (!Xd_0__inst_mult_11_31_q  $ (((Xd_0__inst_mult_11_28_q  & Xd_0__inst_mult_11_29_q )))) ) + ( Xd_0__inst_mult_11_234  ) + ( Xd_0__inst_mult_11_233  ))
// Xd_0__inst_mult_11_237  = CARRY(( !Xd_0__inst_mult_11_30_q  $ (!Xd_0__inst_mult_11_31_q  $ (((Xd_0__inst_mult_11_28_q  & Xd_0__inst_mult_11_29_q )))) ) + ( Xd_0__inst_mult_11_234  ) + ( Xd_0__inst_mult_11_233  ))
// Xd_0__inst_mult_11_238  = SHARE((Xd_0__inst_mult_11_28_q  & (Xd_0__inst_mult_11_29_q  & (!Xd_0__inst_mult_11_30_q  $ (!Xd_0__inst_mult_11_31_q )))))

	.dataa(!Xd_0__inst_mult_11_30_q ),
	.datab(!Xd_0__inst_mult_11_31_q ),
	.datac(!Xd_0__inst_mult_11_28_q ),
	.datad(!Xd_0__inst_mult_11_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_233 ),
	.sharein(Xd_0__inst_mult_11_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_236 ),
	.cout(Xd_0__inst_mult_11_237 ),
	.shareout(Xd_0__inst_mult_11_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_84 (
// Equation(s):
// Xd_0__inst_mult_8_236  = SUM(( !Xd_0__inst_mult_8_30_q  $ (!Xd_0__inst_mult_8_31_q  $ (((Xd_0__inst_mult_8_28_q  & Xd_0__inst_mult_8_29_q )))) ) + ( Xd_0__inst_mult_8_234  ) + ( Xd_0__inst_mult_8_233  ))
// Xd_0__inst_mult_8_237  = CARRY(( !Xd_0__inst_mult_8_30_q  $ (!Xd_0__inst_mult_8_31_q  $ (((Xd_0__inst_mult_8_28_q  & Xd_0__inst_mult_8_29_q )))) ) + ( Xd_0__inst_mult_8_234  ) + ( Xd_0__inst_mult_8_233  ))
// Xd_0__inst_mult_8_238  = SHARE((Xd_0__inst_mult_8_28_q  & (Xd_0__inst_mult_8_29_q  & (!Xd_0__inst_mult_8_30_q  $ (!Xd_0__inst_mult_8_31_q )))))

	.dataa(!Xd_0__inst_mult_8_30_q ),
	.datab(!Xd_0__inst_mult_8_31_q ),
	.datac(!Xd_0__inst_mult_8_28_q ),
	.datad(!Xd_0__inst_mult_8_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_233 ),
	.sharein(Xd_0__inst_mult_8_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_236 ),
	.cout(Xd_0__inst_mult_8_237 ),
	.shareout(Xd_0__inst_mult_8_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_80 (
// Equation(s):
// Xd_0__inst_mult_9_232  = SUM(( !Xd_0__inst_mult_9_30_q  $ (!Xd_0__inst_mult_9_31_q  $ (((Xd_0__inst_mult_9_28_q  & Xd_0__inst_mult_9_29_q )))) ) + ( Xd_0__inst_mult_9_230  ) + ( Xd_0__inst_mult_9_229  ))
// Xd_0__inst_mult_9_233  = CARRY(( !Xd_0__inst_mult_9_30_q  $ (!Xd_0__inst_mult_9_31_q  $ (((Xd_0__inst_mult_9_28_q  & Xd_0__inst_mult_9_29_q )))) ) + ( Xd_0__inst_mult_9_230  ) + ( Xd_0__inst_mult_9_229  ))
// Xd_0__inst_mult_9_234  = SHARE((Xd_0__inst_mult_9_28_q  & (Xd_0__inst_mult_9_29_q  & (!Xd_0__inst_mult_9_30_q  $ (!Xd_0__inst_mult_9_31_q )))))

	.dataa(!Xd_0__inst_mult_9_30_q ),
	.datab(!Xd_0__inst_mult_9_31_q ),
	.datac(!Xd_0__inst_mult_9_28_q ),
	.datad(!Xd_0__inst_mult_9_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_229 ),
	.sharein(Xd_0__inst_mult_9_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_232 ),
	.cout(Xd_0__inst_mult_9_233 ),
	.shareout(Xd_0__inst_mult_9_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_80 (
// Equation(s):
// Xd_0__inst_mult_6_232  = SUM(( !Xd_0__inst_mult_6_30_q  $ (!Xd_0__inst_mult_6_31_q  $ (((Xd_0__inst_mult_6_28_q  & Xd_0__inst_mult_6_29_q )))) ) + ( Xd_0__inst_mult_6_230  ) + ( Xd_0__inst_mult_6_229  ))
// Xd_0__inst_mult_6_233  = CARRY(( !Xd_0__inst_mult_6_30_q  $ (!Xd_0__inst_mult_6_31_q  $ (((Xd_0__inst_mult_6_28_q  & Xd_0__inst_mult_6_29_q )))) ) + ( Xd_0__inst_mult_6_230  ) + ( Xd_0__inst_mult_6_229  ))
// Xd_0__inst_mult_6_234  = SHARE((Xd_0__inst_mult_6_28_q  & (Xd_0__inst_mult_6_29_q  & (!Xd_0__inst_mult_6_30_q  $ (!Xd_0__inst_mult_6_31_q )))))

	.dataa(!Xd_0__inst_mult_6_30_q ),
	.datab(!Xd_0__inst_mult_6_31_q ),
	.datac(!Xd_0__inst_mult_6_28_q ),
	.datad(!Xd_0__inst_mult_6_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_229 ),
	.sharein(Xd_0__inst_mult_6_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_232 ),
	.cout(Xd_0__inst_mult_6_233 ),
	.shareout(Xd_0__inst_mult_6_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_78 (
// Equation(s):
// Xd_0__inst_mult_7_224  = SUM(( !Xd_0__inst_mult_7_30_q  $ (!Xd_0__inst_mult_7_31_q  $ (((Xd_0__inst_mult_7_28_q  & Xd_0__inst_mult_7_29_q )))) ) + ( Xd_0__inst_mult_7_222  ) + ( Xd_0__inst_mult_7_221  ))
// Xd_0__inst_mult_7_225  = CARRY(( !Xd_0__inst_mult_7_30_q  $ (!Xd_0__inst_mult_7_31_q  $ (((Xd_0__inst_mult_7_28_q  & Xd_0__inst_mult_7_29_q )))) ) + ( Xd_0__inst_mult_7_222  ) + ( Xd_0__inst_mult_7_221  ))
// Xd_0__inst_mult_7_226  = SHARE((Xd_0__inst_mult_7_28_q  & (Xd_0__inst_mult_7_29_q  & (!Xd_0__inst_mult_7_30_q  $ (!Xd_0__inst_mult_7_31_q )))))

	.dataa(!Xd_0__inst_mult_7_30_q ),
	.datab(!Xd_0__inst_mult_7_31_q ),
	.datac(!Xd_0__inst_mult_7_28_q ),
	.datad(!Xd_0__inst_mult_7_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_221 ),
	.sharein(Xd_0__inst_mult_7_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_224 ),
	.cout(Xd_0__inst_mult_7_225 ),
	.shareout(Xd_0__inst_mult_7_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_88 (
// Equation(s):
// Xd_0__inst_mult_4_252  = SUM(( !Xd_0__inst_mult_4_30_q  $ (!Xd_0__inst_mult_4_31_q  $ (((Xd_0__inst_mult_4_28_q  & Xd_0__inst_mult_4_29_q )))) ) + ( Xd_0__inst_mult_4_250  ) + ( Xd_0__inst_mult_4_249  ))
// Xd_0__inst_mult_4_253  = CARRY(( !Xd_0__inst_mult_4_30_q  $ (!Xd_0__inst_mult_4_31_q  $ (((Xd_0__inst_mult_4_28_q  & Xd_0__inst_mult_4_29_q )))) ) + ( Xd_0__inst_mult_4_250  ) + ( Xd_0__inst_mult_4_249  ))
// Xd_0__inst_mult_4_254  = SHARE((Xd_0__inst_mult_4_28_q  & (Xd_0__inst_mult_4_29_q  & (!Xd_0__inst_mult_4_30_q  $ (!Xd_0__inst_mult_4_31_q )))))

	.dataa(!Xd_0__inst_mult_4_30_q ),
	.datab(!Xd_0__inst_mult_4_31_q ),
	.datac(!Xd_0__inst_mult_4_28_q ),
	.datad(!Xd_0__inst_mult_4_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_249 ),
	.sharein(Xd_0__inst_mult_4_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_252 ),
	.cout(Xd_0__inst_mult_4_253 ),
	.shareout(Xd_0__inst_mult_4_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_78 (
// Equation(s):
// Xd_0__inst_mult_5_224  = SUM(( !Xd_0__inst_mult_5_30_q  $ (!Xd_0__inst_mult_5_31_q  $ (((Xd_0__inst_mult_5_28_q  & Xd_0__inst_mult_5_29_q )))) ) + ( Xd_0__inst_mult_5_222  ) + ( Xd_0__inst_mult_5_221  ))
// Xd_0__inst_mult_5_225  = CARRY(( !Xd_0__inst_mult_5_30_q  $ (!Xd_0__inst_mult_5_31_q  $ (((Xd_0__inst_mult_5_28_q  & Xd_0__inst_mult_5_29_q )))) ) + ( Xd_0__inst_mult_5_222  ) + ( Xd_0__inst_mult_5_221  ))
// Xd_0__inst_mult_5_226  = SHARE((Xd_0__inst_mult_5_28_q  & (Xd_0__inst_mult_5_29_q  & (!Xd_0__inst_mult_5_30_q  $ (!Xd_0__inst_mult_5_31_q )))))

	.dataa(!Xd_0__inst_mult_5_30_q ),
	.datab(!Xd_0__inst_mult_5_31_q ),
	.datac(!Xd_0__inst_mult_5_28_q ),
	.datad(!Xd_0__inst_mult_5_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_221 ),
	.sharein(Xd_0__inst_mult_5_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_224 ),
	.cout(Xd_0__inst_mult_5_225 ),
	.shareout(Xd_0__inst_mult_5_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_82 (
// Equation(s):
// Xd_0__inst_mult_2_228  = SUM(( !Xd_0__inst_mult_2_30_q  $ (!Xd_0__inst_mult_2_31_q  $ (((Xd_0__inst_mult_2_28_q  & Xd_0__inst_mult_2_29_q )))) ) + ( Xd_0__inst_mult_2_226  ) + ( Xd_0__inst_mult_2_225  ))
// Xd_0__inst_mult_2_229  = CARRY(( !Xd_0__inst_mult_2_30_q  $ (!Xd_0__inst_mult_2_31_q  $ (((Xd_0__inst_mult_2_28_q  & Xd_0__inst_mult_2_29_q )))) ) + ( Xd_0__inst_mult_2_226  ) + ( Xd_0__inst_mult_2_225  ))
// Xd_0__inst_mult_2_230  = SHARE((Xd_0__inst_mult_2_28_q  & (Xd_0__inst_mult_2_29_q  & (!Xd_0__inst_mult_2_30_q  $ (!Xd_0__inst_mult_2_31_q )))))

	.dataa(!Xd_0__inst_mult_2_30_q ),
	.datab(!Xd_0__inst_mult_2_31_q ),
	.datac(!Xd_0__inst_mult_2_28_q ),
	.datad(!Xd_0__inst_mult_2_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_225 ),
	.sharein(Xd_0__inst_mult_2_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_228 ),
	.cout(Xd_0__inst_mult_2_229 ),
	.shareout(Xd_0__inst_mult_2_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_78 (
// Equation(s):
// Xd_0__inst_mult_3_224  = SUM(( !Xd_0__inst_mult_3_30_q  $ (!Xd_0__inst_mult_3_31_q  $ (((Xd_0__inst_mult_3_28_q  & Xd_0__inst_mult_3_29_q )))) ) + ( Xd_0__inst_mult_3_222  ) + ( Xd_0__inst_mult_3_221  ))
// Xd_0__inst_mult_3_225  = CARRY(( !Xd_0__inst_mult_3_30_q  $ (!Xd_0__inst_mult_3_31_q  $ (((Xd_0__inst_mult_3_28_q  & Xd_0__inst_mult_3_29_q )))) ) + ( Xd_0__inst_mult_3_222  ) + ( Xd_0__inst_mult_3_221  ))
// Xd_0__inst_mult_3_226  = SHARE((Xd_0__inst_mult_3_28_q  & (Xd_0__inst_mult_3_29_q  & (!Xd_0__inst_mult_3_30_q  $ (!Xd_0__inst_mult_3_31_q )))))

	.dataa(!Xd_0__inst_mult_3_30_q ),
	.datab(!Xd_0__inst_mult_3_31_q ),
	.datac(!Xd_0__inst_mult_3_28_q ),
	.datad(!Xd_0__inst_mult_3_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_221 ),
	.sharein(Xd_0__inst_mult_3_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_224 ),
	.cout(Xd_0__inst_mult_3_225 ),
	.shareout(Xd_0__inst_mult_3_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_82 (
// Equation(s):
// Xd_0__inst_mult_0_228  = SUM(( !Xd_0__inst_mult_0_30_q  $ (!Xd_0__inst_mult_0_31_q  $ (((Xd_0__inst_mult_0_28_q  & Xd_0__inst_mult_0_29_q )))) ) + ( Xd_0__inst_mult_0_226  ) + ( Xd_0__inst_mult_0_225  ))
// Xd_0__inst_mult_0_229  = CARRY(( !Xd_0__inst_mult_0_30_q  $ (!Xd_0__inst_mult_0_31_q  $ (((Xd_0__inst_mult_0_28_q  & Xd_0__inst_mult_0_29_q )))) ) + ( Xd_0__inst_mult_0_226  ) + ( Xd_0__inst_mult_0_225  ))
// Xd_0__inst_mult_0_230  = SHARE((Xd_0__inst_mult_0_28_q  & (Xd_0__inst_mult_0_29_q  & (!Xd_0__inst_mult_0_30_q  $ (!Xd_0__inst_mult_0_31_q )))))

	.dataa(!Xd_0__inst_mult_0_30_q ),
	.datab(!Xd_0__inst_mult_0_31_q ),
	.datac(!Xd_0__inst_mult_0_28_q ),
	.datad(!Xd_0__inst_mult_0_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_225 ),
	.sharein(Xd_0__inst_mult_0_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_228 ),
	.cout(Xd_0__inst_mult_0_229 ),
	.shareout(Xd_0__inst_mult_0_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_82 (
// Equation(s):
// Xd_0__inst_mult_1_228  = SUM(( !Xd_0__inst_mult_1_30_q  $ (!Xd_0__inst_mult_1_31_q  $ (((Xd_0__inst_mult_1_28_q  & Xd_0__inst_mult_1_29_q )))) ) + ( Xd_0__inst_mult_1_226  ) + ( Xd_0__inst_mult_1_225  ))
// Xd_0__inst_mult_1_229  = CARRY(( !Xd_0__inst_mult_1_30_q  $ (!Xd_0__inst_mult_1_31_q  $ (((Xd_0__inst_mult_1_28_q  & Xd_0__inst_mult_1_29_q )))) ) + ( Xd_0__inst_mult_1_226  ) + ( Xd_0__inst_mult_1_225  ))
// Xd_0__inst_mult_1_230  = SHARE((Xd_0__inst_mult_1_28_q  & (Xd_0__inst_mult_1_29_q  & (!Xd_0__inst_mult_1_30_q  $ (!Xd_0__inst_mult_1_31_q )))))

	.dataa(!Xd_0__inst_mult_1_30_q ),
	.datab(!Xd_0__inst_mult_1_31_q ),
	.datac(!Xd_0__inst_mult_1_28_q ),
	.datad(!Xd_0__inst_mult_1_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_225 ),
	.sharein(Xd_0__inst_mult_1_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_228 ),
	.cout(Xd_0__inst_mult_1_229 ),
	.shareout(Xd_0__inst_mult_1_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_85 (
// Equation(s):
// Xd_0__inst_mult_12_252  = SUM(( !Xd_0__inst_mult_12_32_q  $ (!Xd_0__inst_mult_12_33_q  $ (((Xd_0__inst_mult_12_30_q  & Xd_0__inst_mult_12_31_q )))) ) + ( Xd_0__inst_mult_12_250  ) + ( Xd_0__inst_mult_12_249  ))
// Xd_0__inst_mult_12_253  = CARRY(( !Xd_0__inst_mult_12_32_q  $ (!Xd_0__inst_mult_12_33_q  $ (((Xd_0__inst_mult_12_30_q  & Xd_0__inst_mult_12_31_q )))) ) + ( Xd_0__inst_mult_12_250  ) + ( Xd_0__inst_mult_12_249  ))
// Xd_0__inst_mult_12_254  = SHARE((Xd_0__inst_mult_12_30_q  & (Xd_0__inst_mult_12_31_q  & (!Xd_0__inst_mult_12_32_q  $ (!Xd_0__inst_mult_12_33_q )))))

	.dataa(!Xd_0__inst_mult_12_32_q ),
	.datab(!Xd_0__inst_mult_12_33_q ),
	.datac(!Xd_0__inst_mult_12_30_q ),
	.datad(!Xd_0__inst_mult_12_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_249 ),
	.sharein(Xd_0__inst_mult_12_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_252 ),
	.cout(Xd_0__inst_mult_12_253 ),
	.shareout(Xd_0__inst_mult_12_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_85 (
// Equation(s):
// Xd_0__inst_mult_13_240  = SUM(( !Xd_0__inst_mult_13_32_q  $ (!Xd_0__inst_mult_13_33_q  $ (((Xd_0__inst_mult_13_30_q  & Xd_0__inst_mult_13_31_q )))) ) + ( Xd_0__inst_mult_13_238  ) + ( Xd_0__inst_mult_13_237  ))
// Xd_0__inst_mult_13_241  = CARRY(( !Xd_0__inst_mult_13_32_q  $ (!Xd_0__inst_mult_13_33_q  $ (((Xd_0__inst_mult_13_30_q  & Xd_0__inst_mult_13_31_q )))) ) + ( Xd_0__inst_mult_13_238  ) + ( Xd_0__inst_mult_13_237  ))
// Xd_0__inst_mult_13_242  = SHARE((Xd_0__inst_mult_13_30_q  & (Xd_0__inst_mult_13_31_q  & (!Xd_0__inst_mult_13_32_q  $ (!Xd_0__inst_mult_13_33_q )))))

	.dataa(!Xd_0__inst_mult_13_32_q ),
	.datab(!Xd_0__inst_mult_13_33_q ),
	.datac(!Xd_0__inst_mult_13_30_q ),
	.datad(!Xd_0__inst_mult_13_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_237 ),
	.sharein(Xd_0__inst_mult_13_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_240 ),
	.cout(Xd_0__inst_mult_13_241 ),
	.shareout(Xd_0__inst_mult_13_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_89 (
// Equation(s):
// Xd_0__inst_mult_14_256  = SUM(( !Xd_0__inst_mult_14_32_q  $ (!Xd_0__inst_mult_14_33_q  $ (((Xd_0__inst_mult_14_30_q  & Xd_0__inst_mult_14_31_q )))) ) + ( Xd_0__inst_mult_14_254  ) + ( Xd_0__inst_mult_14_253  ))
// Xd_0__inst_mult_14_257  = CARRY(( !Xd_0__inst_mult_14_32_q  $ (!Xd_0__inst_mult_14_33_q  $ (((Xd_0__inst_mult_14_30_q  & Xd_0__inst_mult_14_31_q )))) ) + ( Xd_0__inst_mult_14_254  ) + ( Xd_0__inst_mult_14_253  ))
// Xd_0__inst_mult_14_258  = SHARE((Xd_0__inst_mult_14_30_q  & (Xd_0__inst_mult_14_31_q  & (!Xd_0__inst_mult_14_32_q  $ (!Xd_0__inst_mult_14_33_q )))))

	.dataa(!Xd_0__inst_mult_14_32_q ),
	.datab(!Xd_0__inst_mult_14_33_q ),
	.datac(!Xd_0__inst_mult_14_30_q ),
	.datad(!Xd_0__inst_mult_14_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_253 ),
	.sharein(Xd_0__inst_mult_14_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_256 ),
	.cout(Xd_0__inst_mult_14_257 ),
	.shareout(Xd_0__inst_mult_14_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_89 (
// Equation(s):
// Xd_0__inst_mult_15_256  = SUM(( !Xd_0__inst_mult_15_32_q  $ (!Xd_0__inst_mult_15_33_q  $ (((Xd_0__inst_mult_15_30_q  & Xd_0__inst_mult_15_31_q )))) ) + ( Xd_0__inst_mult_15_254  ) + ( Xd_0__inst_mult_15_253  ))
// Xd_0__inst_mult_15_257  = CARRY(( !Xd_0__inst_mult_15_32_q  $ (!Xd_0__inst_mult_15_33_q  $ (((Xd_0__inst_mult_15_30_q  & Xd_0__inst_mult_15_31_q )))) ) + ( Xd_0__inst_mult_15_254  ) + ( Xd_0__inst_mult_15_253  ))
// Xd_0__inst_mult_15_258  = SHARE((Xd_0__inst_mult_15_30_q  & (Xd_0__inst_mult_15_31_q  & (!Xd_0__inst_mult_15_32_q  $ (!Xd_0__inst_mult_15_33_q )))))

	.dataa(!Xd_0__inst_mult_15_32_q ),
	.datab(!Xd_0__inst_mult_15_33_q ),
	.datac(!Xd_0__inst_mult_15_30_q ),
	.datad(!Xd_0__inst_mult_15_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_253 ),
	.sharein(Xd_0__inst_mult_15_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_256 ),
	.cout(Xd_0__inst_mult_15_257 ),
	.shareout(Xd_0__inst_mult_15_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_81 (
// Equation(s):
// Xd_0__inst_mult_10_236  = SUM(( !Xd_0__inst_mult_10_32_q  $ (!Xd_0__inst_mult_10_33_q  $ (((Xd_0__inst_mult_10_30_q  & Xd_0__inst_mult_10_31_q )))) ) + ( Xd_0__inst_mult_10_234  ) + ( Xd_0__inst_mult_10_233  ))
// Xd_0__inst_mult_10_237  = CARRY(( !Xd_0__inst_mult_10_32_q  $ (!Xd_0__inst_mult_10_33_q  $ (((Xd_0__inst_mult_10_30_q  & Xd_0__inst_mult_10_31_q )))) ) + ( Xd_0__inst_mult_10_234  ) + ( Xd_0__inst_mult_10_233  ))
// Xd_0__inst_mult_10_238  = SHARE((Xd_0__inst_mult_10_30_q  & (Xd_0__inst_mult_10_31_q  & (!Xd_0__inst_mult_10_32_q  $ (!Xd_0__inst_mult_10_33_q )))))

	.dataa(!Xd_0__inst_mult_10_32_q ),
	.datab(!Xd_0__inst_mult_10_33_q ),
	.datac(!Xd_0__inst_mult_10_30_q ),
	.datad(!Xd_0__inst_mult_10_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_233 ),
	.sharein(Xd_0__inst_mult_10_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_236 ),
	.cout(Xd_0__inst_mult_10_237 ),
	.shareout(Xd_0__inst_mult_10_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_85 (
// Equation(s):
// Xd_0__inst_mult_11_240  = SUM(( !Xd_0__inst_mult_11_32_q  $ (!Xd_0__inst_mult_11_33_q  $ (((Xd_0__inst_mult_11_30_q  & Xd_0__inst_mult_11_31_q )))) ) + ( Xd_0__inst_mult_11_238  ) + ( Xd_0__inst_mult_11_237  ))
// Xd_0__inst_mult_11_241  = CARRY(( !Xd_0__inst_mult_11_32_q  $ (!Xd_0__inst_mult_11_33_q  $ (((Xd_0__inst_mult_11_30_q  & Xd_0__inst_mult_11_31_q )))) ) + ( Xd_0__inst_mult_11_238  ) + ( Xd_0__inst_mult_11_237  ))
// Xd_0__inst_mult_11_242  = SHARE((Xd_0__inst_mult_11_30_q  & (Xd_0__inst_mult_11_31_q  & (!Xd_0__inst_mult_11_32_q  $ (!Xd_0__inst_mult_11_33_q )))))

	.dataa(!Xd_0__inst_mult_11_32_q ),
	.datab(!Xd_0__inst_mult_11_33_q ),
	.datac(!Xd_0__inst_mult_11_30_q ),
	.datad(!Xd_0__inst_mult_11_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_237 ),
	.sharein(Xd_0__inst_mult_11_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_240 ),
	.cout(Xd_0__inst_mult_11_241 ),
	.shareout(Xd_0__inst_mult_11_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_85 (
// Equation(s):
// Xd_0__inst_mult_8_240  = SUM(( !Xd_0__inst_mult_8_32_q  $ (!Xd_0__inst_mult_8_33_q  $ (((Xd_0__inst_mult_8_30_q  & Xd_0__inst_mult_8_31_q )))) ) + ( Xd_0__inst_mult_8_238  ) + ( Xd_0__inst_mult_8_237  ))
// Xd_0__inst_mult_8_241  = CARRY(( !Xd_0__inst_mult_8_32_q  $ (!Xd_0__inst_mult_8_33_q  $ (((Xd_0__inst_mult_8_30_q  & Xd_0__inst_mult_8_31_q )))) ) + ( Xd_0__inst_mult_8_238  ) + ( Xd_0__inst_mult_8_237  ))
// Xd_0__inst_mult_8_242  = SHARE((Xd_0__inst_mult_8_30_q  & (Xd_0__inst_mult_8_31_q  & (!Xd_0__inst_mult_8_32_q  $ (!Xd_0__inst_mult_8_33_q )))))

	.dataa(!Xd_0__inst_mult_8_32_q ),
	.datab(!Xd_0__inst_mult_8_33_q ),
	.datac(!Xd_0__inst_mult_8_30_q ),
	.datad(!Xd_0__inst_mult_8_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_237 ),
	.sharein(Xd_0__inst_mult_8_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_240 ),
	.cout(Xd_0__inst_mult_8_241 ),
	.shareout(Xd_0__inst_mult_8_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_81 (
// Equation(s):
// Xd_0__inst_mult_9_236  = SUM(( !Xd_0__inst_mult_9_32_q  $ (!Xd_0__inst_mult_9_33_q  $ (((Xd_0__inst_mult_9_30_q  & Xd_0__inst_mult_9_31_q )))) ) + ( Xd_0__inst_mult_9_234  ) + ( Xd_0__inst_mult_9_233  ))
// Xd_0__inst_mult_9_237  = CARRY(( !Xd_0__inst_mult_9_32_q  $ (!Xd_0__inst_mult_9_33_q  $ (((Xd_0__inst_mult_9_30_q  & Xd_0__inst_mult_9_31_q )))) ) + ( Xd_0__inst_mult_9_234  ) + ( Xd_0__inst_mult_9_233  ))
// Xd_0__inst_mult_9_238  = SHARE((Xd_0__inst_mult_9_30_q  & (Xd_0__inst_mult_9_31_q  & (!Xd_0__inst_mult_9_32_q  $ (!Xd_0__inst_mult_9_33_q )))))

	.dataa(!Xd_0__inst_mult_9_32_q ),
	.datab(!Xd_0__inst_mult_9_33_q ),
	.datac(!Xd_0__inst_mult_9_30_q ),
	.datad(!Xd_0__inst_mult_9_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_233 ),
	.sharein(Xd_0__inst_mult_9_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_236 ),
	.cout(Xd_0__inst_mult_9_237 ),
	.shareout(Xd_0__inst_mult_9_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_81 (
// Equation(s):
// Xd_0__inst_mult_6_236  = SUM(( !Xd_0__inst_mult_6_32_q  $ (!Xd_0__inst_mult_6_33_q  $ (((Xd_0__inst_mult_6_30_q  & Xd_0__inst_mult_6_31_q )))) ) + ( Xd_0__inst_mult_6_234  ) + ( Xd_0__inst_mult_6_233  ))
// Xd_0__inst_mult_6_237  = CARRY(( !Xd_0__inst_mult_6_32_q  $ (!Xd_0__inst_mult_6_33_q  $ (((Xd_0__inst_mult_6_30_q  & Xd_0__inst_mult_6_31_q )))) ) + ( Xd_0__inst_mult_6_234  ) + ( Xd_0__inst_mult_6_233  ))
// Xd_0__inst_mult_6_238  = SHARE((Xd_0__inst_mult_6_30_q  & (Xd_0__inst_mult_6_31_q  & (!Xd_0__inst_mult_6_32_q  $ (!Xd_0__inst_mult_6_33_q )))))

	.dataa(!Xd_0__inst_mult_6_32_q ),
	.datab(!Xd_0__inst_mult_6_33_q ),
	.datac(!Xd_0__inst_mult_6_30_q ),
	.datad(!Xd_0__inst_mult_6_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_233 ),
	.sharein(Xd_0__inst_mult_6_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_236 ),
	.cout(Xd_0__inst_mult_6_237 ),
	.shareout(Xd_0__inst_mult_6_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_79 (
// Equation(s):
// Xd_0__inst_mult_7_228  = SUM(( !Xd_0__inst_mult_7_32_q  $ (!Xd_0__inst_mult_7_33_q  $ (((Xd_0__inst_mult_7_30_q  & Xd_0__inst_mult_7_31_q )))) ) + ( Xd_0__inst_mult_7_226  ) + ( Xd_0__inst_mult_7_225  ))
// Xd_0__inst_mult_7_229  = CARRY(( !Xd_0__inst_mult_7_32_q  $ (!Xd_0__inst_mult_7_33_q  $ (((Xd_0__inst_mult_7_30_q  & Xd_0__inst_mult_7_31_q )))) ) + ( Xd_0__inst_mult_7_226  ) + ( Xd_0__inst_mult_7_225  ))
// Xd_0__inst_mult_7_230  = SHARE((Xd_0__inst_mult_7_30_q  & (Xd_0__inst_mult_7_31_q  & (!Xd_0__inst_mult_7_32_q  $ (!Xd_0__inst_mult_7_33_q )))))

	.dataa(!Xd_0__inst_mult_7_32_q ),
	.datab(!Xd_0__inst_mult_7_33_q ),
	.datac(!Xd_0__inst_mult_7_30_q ),
	.datad(!Xd_0__inst_mult_7_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_225 ),
	.sharein(Xd_0__inst_mult_7_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_228 ),
	.cout(Xd_0__inst_mult_7_229 ),
	.shareout(Xd_0__inst_mult_7_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_89 (
// Equation(s):
// Xd_0__inst_mult_4_256  = SUM(( !Xd_0__inst_mult_4_32_q  $ (!Xd_0__inst_mult_4_33_q  $ (((Xd_0__inst_mult_4_30_q  & Xd_0__inst_mult_4_31_q )))) ) + ( Xd_0__inst_mult_4_254  ) + ( Xd_0__inst_mult_4_253  ))
// Xd_0__inst_mult_4_257  = CARRY(( !Xd_0__inst_mult_4_32_q  $ (!Xd_0__inst_mult_4_33_q  $ (((Xd_0__inst_mult_4_30_q  & Xd_0__inst_mult_4_31_q )))) ) + ( Xd_0__inst_mult_4_254  ) + ( Xd_0__inst_mult_4_253  ))
// Xd_0__inst_mult_4_258  = SHARE((Xd_0__inst_mult_4_30_q  & (Xd_0__inst_mult_4_31_q  & (!Xd_0__inst_mult_4_32_q  $ (!Xd_0__inst_mult_4_33_q )))))

	.dataa(!Xd_0__inst_mult_4_32_q ),
	.datab(!Xd_0__inst_mult_4_33_q ),
	.datac(!Xd_0__inst_mult_4_30_q ),
	.datad(!Xd_0__inst_mult_4_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_253 ),
	.sharein(Xd_0__inst_mult_4_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_256 ),
	.cout(Xd_0__inst_mult_4_257 ),
	.shareout(Xd_0__inst_mult_4_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_79 (
// Equation(s):
// Xd_0__inst_mult_5_228  = SUM(( !Xd_0__inst_mult_5_32_q  $ (!Xd_0__inst_mult_5_33_q  $ (((Xd_0__inst_mult_5_30_q  & Xd_0__inst_mult_5_31_q )))) ) + ( Xd_0__inst_mult_5_226  ) + ( Xd_0__inst_mult_5_225  ))
// Xd_0__inst_mult_5_229  = CARRY(( !Xd_0__inst_mult_5_32_q  $ (!Xd_0__inst_mult_5_33_q  $ (((Xd_0__inst_mult_5_30_q  & Xd_0__inst_mult_5_31_q )))) ) + ( Xd_0__inst_mult_5_226  ) + ( Xd_0__inst_mult_5_225  ))
// Xd_0__inst_mult_5_230  = SHARE((Xd_0__inst_mult_5_30_q  & (Xd_0__inst_mult_5_31_q  & (!Xd_0__inst_mult_5_32_q  $ (!Xd_0__inst_mult_5_33_q )))))

	.dataa(!Xd_0__inst_mult_5_32_q ),
	.datab(!Xd_0__inst_mult_5_33_q ),
	.datac(!Xd_0__inst_mult_5_30_q ),
	.datad(!Xd_0__inst_mult_5_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_225 ),
	.sharein(Xd_0__inst_mult_5_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_228 ),
	.cout(Xd_0__inst_mult_5_229 ),
	.shareout(Xd_0__inst_mult_5_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_83 (
// Equation(s):
// Xd_0__inst_mult_2_232  = SUM(( !Xd_0__inst_mult_2_32_q  $ (!Xd_0__inst_mult_2_33_q  $ (((Xd_0__inst_mult_2_30_q  & Xd_0__inst_mult_2_31_q )))) ) + ( Xd_0__inst_mult_2_230  ) + ( Xd_0__inst_mult_2_229  ))
// Xd_0__inst_mult_2_233  = CARRY(( !Xd_0__inst_mult_2_32_q  $ (!Xd_0__inst_mult_2_33_q  $ (((Xd_0__inst_mult_2_30_q  & Xd_0__inst_mult_2_31_q )))) ) + ( Xd_0__inst_mult_2_230  ) + ( Xd_0__inst_mult_2_229  ))
// Xd_0__inst_mult_2_234  = SHARE((Xd_0__inst_mult_2_30_q  & (Xd_0__inst_mult_2_31_q  & (!Xd_0__inst_mult_2_32_q  $ (!Xd_0__inst_mult_2_33_q )))))

	.dataa(!Xd_0__inst_mult_2_32_q ),
	.datab(!Xd_0__inst_mult_2_33_q ),
	.datac(!Xd_0__inst_mult_2_30_q ),
	.datad(!Xd_0__inst_mult_2_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_229 ),
	.sharein(Xd_0__inst_mult_2_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_232 ),
	.cout(Xd_0__inst_mult_2_233 ),
	.shareout(Xd_0__inst_mult_2_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_79 (
// Equation(s):
// Xd_0__inst_mult_3_228  = SUM(( !Xd_0__inst_mult_3_32_q  $ (!Xd_0__inst_mult_3_33_q  $ (((Xd_0__inst_mult_3_30_q  & Xd_0__inst_mult_3_31_q )))) ) + ( Xd_0__inst_mult_3_226  ) + ( Xd_0__inst_mult_3_225  ))
// Xd_0__inst_mult_3_229  = CARRY(( !Xd_0__inst_mult_3_32_q  $ (!Xd_0__inst_mult_3_33_q  $ (((Xd_0__inst_mult_3_30_q  & Xd_0__inst_mult_3_31_q )))) ) + ( Xd_0__inst_mult_3_226  ) + ( Xd_0__inst_mult_3_225  ))
// Xd_0__inst_mult_3_230  = SHARE((Xd_0__inst_mult_3_30_q  & (Xd_0__inst_mult_3_31_q  & (!Xd_0__inst_mult_3_32_q  $ (!Xd_0__inst_mult_3_33_q )))))

	.dataa(!Xd_0__inst_mult_3_32_q ),
	.datab(!Xd_0__inst_mult_3_33_q ),
	.datac(!Xd_0__inst_mult_3_30_q ),
	.datad(!Xd_0__inst_mult_3_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_225 ),
	.sharein(Xd_0__inst_mult_3_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_228 ),
	.cout(Xd_0__inst_mult_3_229 ),
	.shareout(Xd_0__inst_mult_3_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_83 (
// Equation(s):
// Xd_0__inst_mult_0_232  = SUM(( !Xd_0__inst_mult_0_32_q  $ (!Xd_0__inst_mult_0_33_q  $ (((Xd_0__inst_mult_0_30_q  & Xd_0__inst_mult_0_31_q )))) ) + ( Xd_0__inst_mult_0_230  ) + ( Xd_0__inst_mult_0_229  ))
// Xd_0__inst_mult_0_233  = CARRY(( !Xd_0__inst_mult_0_32_q  $ (!Xd_0__inst_mult_0_33_q  $ (((Xd_0__inst_mult_0_30_q  & Xd_0__inst_mult_0_31_q )))) ) + ( Xd_0__inst_mult_0_230  ) + ( Xd_0__inst_mult_0_229  ))
// Xd_0__inst_mult_0_234  = SHARE((Xd_0__inst_mult_0_30_q  & (Xd_0__inst_mult_0_31_q  & (!Xd_0__inst_mult_0_32_q  $ (!Xd_0__inst_mult_0_33_q )))))

	.dataa(!Xd_0__inst_mult_0_32_q ),
	.datab(!Xd_0__inst_mult_0_33_q ),
	.datac(!Xd_0__inst_mult_0_30_q ),
	.datad(!Xd_0__inst_mult_0_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_229 ),
	.sharein(Xd_0__inst_mult_0_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_232 ),
	.cout(Xd_0__inst_mult_0_233 ),
	.shareout(Xd_0__inst_mult_0_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_83 (
// Equation(s):
// Xd_0__inst_mult_1_232  = SUM(( !Xd_0__inst_mult_1_32_q  $ (!Xd_0__inst_mult_1_33_q  $ (((Xd_0__inst_mult_1_30_q  & Xd_0__inst_mult_1_31_q )))) ) + ( Xd_0__inst_mult_1_230  ) + ( Xd_0__inst_mult_1_229  ))
// Xd_0__inst_mult_1_233  = CARRY(( !Xd_0__inst_mult_1_32_q  $ (!Xd_0__inst_mult_1_33_q  $ (((Xd_0__inst_mult_1_30_q  & Xd_0__inst_mult_1_31_q )))) ) + ( Xd_0__inst_mult_1_230  ) + ( Xd_0__inst_mult_1_229  ))
// Xd_0__inst_mult_1_234  = SHARE((Xd_0__inst_mult_1_30_q  & (Xd_0__inst_mult_1_31_q  & (!Xd_0__inst_mult_1_32_q  $ (!Xd_0__inst_mult_1_33_q )))))

	.dataa(!Xd_0__inst_mult_1_32_q ),
	.datab(!Xd_0__inst_mult_1_33_q ),
	.datac(!Xd_0__inst_mult_1_30_q ),
	.datad(!Xd_0__inst_mult_1_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_229 ),
	.sharein(Xd_0__inst_mult_1_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_232 ),
	.cout(Xd_0__inst_mult_1_233 ),
	.shareout(Xd_0__inst_mult_1_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_86 (
// Equation(s):
// Xd_0__inst_mult_12_256  = SUM(( (Xd_0__inst_mult_12_32_q  & Xd_0__inst_mult_12_33_q ) ) + ( Xd_0__inst_mult_12_254  ) + ( Xd_0__inst_mult_12_253  ))

	.dataa(!Xd_0__inst_mult_12_32_q ),
	.datab(!Xd_0__inst_mult_12_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_253 ),
	.sharein(Xd_0__inst_mult_12_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_256 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_86 (
// Equation(s):
// Xd_0__inst_mult_13_244  = SUM(( (Xd_0__inst_mult_13_32_q  & Xd_0__inst_mult_13_33_q ) ) + ( Xd_0__inst_mult_13_242  ) + ( Xd_0__inst_mult_13_241  ))

	.dataa(!Xd_0__inst_mult_13_32_q ),
	.datab(!Xd_0__inst_mult_13_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_241 ),
	.sharein(Xd_0__inst_mult_13_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_244 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_90 (
// Equation(s):
// Xd_0__inst_mult_14_260  = SUM(( (Xd_0__inst_mult_14_32_q  & Xd_0__inst_mult_14_33_q ) ) + ( Xd_0__inst_mult_14_258  ) + ( Xd_0__inst_mult_14_257  ))

	.dataa(!Xd_0__inst_mult_14_32_q ),
	.datab(!Xd_0__inst_mult_14_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_257 ),
	.sharein(Xd_0__inst_mult_14_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_260 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_90 (
// Equation(s):
// Xd_0__inst_mult_15_260  = SUM(( (Xd_0__inst_mult_15_32_q  & Xd_0__inst_mult_15_33_q ) ) + ( Xd_0__inst_mult_15_258  ) + ( Xd_0__inst_mult_15_257  ))

	.dataa(!Xd_0__inst_mult_15_32_q ),
	.datab(!Xd_0__inst_mult_15_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_257 ),
	.sharein(Xd_0__inst_mult_15_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_260 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_82 (
// Equation(s):
// Xd_0__inst_mult_10_240  = SUM(( (Xd_0__inst_mult_10_32_q  & Xd_0__inst_mult_10_33_q ) ) + ( Xd_0__inst_mult_10_238  ) + ( Xd_0__inst_mult_10_237  ))

	.dataa(!Xd_0__inst_mult_10_32_q ),
	.datab(!Xd_0__inst_mult_10_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_237 ),
	.sharein(Xd_0__inst_mult_10_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_240 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_86 (
// Equation(s):
// Xd_0__inst_mult_11_244  = SUM(( (Xd_0__inst_mult_11_32_q  & Xd_0__inst_mult_11_33_q ) ) + ( Xd_0__inst_mult_11_242  ) + ( Xd_0__inst_mult_11_241  ))

	.dataa(!Xd_0__inst_mult_11_32_q ),
	.datab(!Xd_0__inst_mult_11_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_241 ),
	.sharein(Xd_0__inst_mult_11_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_244 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_86 (
// Equation(s):
// Xd_0__inst_mult_8_244  = SUM(( (Xd_0__inst_mult_8_32_q  & Xd_0__inst_mult_8_33_q ) ) + ( Xd_0__inst_mult_8_242  ) + ( Xd_0__inst_mult_8_241  ))

	.dataa(!Xd_0__inst_mult_8_32_q ),
	.datab(!Xd_0__inst_mult_8_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_241 ),
	.sharein(Xd_0__inst_mult_8_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_244 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_82 (
// Equation(s):
// Xd_0__inst_mult_9_240  = SUM(( (Xd_0__inst_mult_9_32_q  & Xd_0__inst_mult_9_33_q ) ) + ( Xd_0__inst_mult_9_238  ) + ( Xd_0__inst_mult_9_237  ))

	.dataa(!Xd_0__inst_mult_9_32_q ),
	.datab(!Xd_0__inst_mult_9_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_237 ),
	.sharein(Xd_0__inst_mult_9_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_240 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_82 (
// Equation(s):
// Xd_0__inst_mult_6_240  = SUM(( (Xd_0__inst_mult_6_32_q  & Xd_0__inst_mult_6_33_q ) ) + ( Xd_0__inst_mult_6_238  ) + ( Xd_0__inst_mult_6_237  ))

	.dataa(!Xd_0__inst_mult_6_32_q ),
	.datab(!Xd_0__inst_mult_6_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_237 ),
	.sharein(Xd_0__inst_mult_6_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_240 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_80 (
// Equation(s):
// Xd_0__inst_mult_7_232  = SUM(( (Xd_0__inst_mult_7_32_q  & Xd_0__inst_mult_7_33_q ) ) + ( Xd_0__inst_mult_7_230  ) + ( Xd_0__inst_mult_7_229  ))

	.dataa(!Xd_0__inst_mult_7_32_q ),
	.datab(!Xd_0__inst_mult_7_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_229 ),
	.sharein(Xd_0__inst_mult_7_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_232 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_90 (
// Equation(s):
// Xd_0__inst_mult_4_260  = SUM(( (Xd_0__inst_mult_4_32_q  & Xd_0__inst_mult_4_33_q ) ) + ( Xd_0__inst_mult_4_258  ) + ( Xd_0__inst_mult_4_257  ))

	.dataa(!Xd_0__inst_mult_4_32_q ),
	.datab(!Xd_0__inst_mult_4_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_257 ),
	.sharein(Xd_0__inst_mult_4_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_260 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_80 (
// Equation(s):
// Xd_0__inst_mult_5_232  = SUM(( (Xd_0__inst_mult_5_32_q  & Xd_0__inst_mult_5_33_q ) ) + ( Xd_0__inst_mult_5_230  ) + ( Xd_0__inst_mult_5_229  ))

	.dataa(!Xd_0__inst_mult_5_32_q ),
	.datab(!Xd_0__inst_mult_5_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_229 ),
	.sharein(Xd_0__inst_mult_5_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_232 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_84 (
// Equation(s):
// Xd_0__inst_mult_2_236  = SUM(( (Xd_0__inst_mult_2_32_q  & Xd_0__inst_mult_2_33_q ) ) + ( Xd_0__inst_mult_2_234  ) + ( Xd_0__inst_mult_2_233  ))

	.dataa(!Xd_0__inst_mult_2_32_q ),
	.datab(!Xd_0__inst_mult_2_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_233 ),
	.sharein(Xd_0__inst_mult_2_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_236 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_80 (
// Equation(s):
// Xd_0__inst_mult_3_232  = SUM(( (Xd_0__inst_mult_3_32_q  & Xd_0__inst_mult_3_33_q ) ) + ( Xd_0__inst_mult_3_230  ) + ( Xd_0__inst_mult_3_229  ))

	.dataa(!Xd_0__inst_mult_3_32_q ),
	.datab(!Xd_0__inst_mult_3_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_229 ),
	.sharein(Xd_0__inst_mult_3_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_232 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_84 (
// Equation(s):
// Xd_0__inst_mult_0_236  = SUM(( (Xd_0__inst_mult_0_32_q  & Xd_0__inst_mult_0_33_q ) ) + ( Xd_0__inst_mult_0_234  ) + ( Xd_0__inst_mult_0_233  ))

	.dataa(!Xd_0__inst_mult_0_32_q ),
	.datab(!Xd_0__inst_mult_0_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_233 ),
	.sharein(Xd_0__inst_mult_0_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_236 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_84 (
// Equation(s):
// Xd_0__inst_mult_1_236  = SUM(( (Xd_0__inst_mult_1_32_q  & Xd_0__inst_mult_1_33_q ) ) + ( Xd_0__inst_mult_1_234  ) + ( Xd_0__inst_mult_1_233  ))

	.dataa(!Xd_0__inst_mult_1_32_q ),
	.datab(!Xd_0__inst_mult_1_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_233 ),
	.sharein(Xd_0__inst_mult_1_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_236 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_87 (
// Equation(s):
// Xd_0__inst_mult_12_260  = SUM(( (din_a[144] & din_b[144]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_261  = CARRY(( (din_a[144] & din_b[144]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_262  = SHARE((din_a[144] & din_b[145]))

	.dataa(!din_a[144]),
	.datab(!din_b[144]),
	.datac(!din_b[145]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_12_260 ),
	.cout(Xd_0__inst_mult_12_261 ),
	.shareout(Xd_0__inst_mult_12_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_87 (
// Equation(s):
// Xd_0__inst_mult_13_248  = SUM(( (din_a[156] & din_b[156]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_249  = CARRY(( (din_a[156] & din_b[156]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_250  = SHARE((din_a[156] & din_b[157]))

	.dataa(!din_a[156]),
	.datab(!din_b[156]),
	.datac(!din_b[157]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_13_248 ),
	.cout(Xd_0__inst_mult_13_249 ),
	.shareout(Xd_0__inst_mult_13_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_1 (
// Equation(s):
// Xd_0__inst_i29_1_sumout  = SUM(( !din_a[155] $ (!din_b[155]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_2  = CARRY(( !din_a[155] $ (!din_b[155]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_3  = SHARE(GND)

	.dataa(!din_a[155]),
	.datab(!din_b[155]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i29_1_sumout ),
	.cout(Xd_0__inst_i29_2 ),
	.shareout(Xd_0__inst_i29_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_5 (
// Equation(s):
// Xd_0__inst_i29_5_sumout  = SUM(( !din_a[167] $ (!din_b[167]) ) + ( Xd_0__inst_i29_3  ) + ( Xd_0__inst_i29_2  ))
// Xd_0__inst_i29_6  = CARRY(( !din_a[167] $ (!din_b[167]) ) + ( Xd_0__inst_i29_3  ) + ( Xd_0__inst_i29_2  ))
// Xd_0__inst_i29_7  = SHARE(GND)

	.dataa(!din_a[167]),
	.datab(!din_b[167]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_2 ),
	.sharein(Xd_0__inst_i29_3 ),
	.combout(),
	.sumout(Xd_0__inst_i29_5_sumout ),
	.cout(Xd_0__inst_i29_6 ),
	.shareout(Xd_0__inst_i29_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_83 (
// Equation(s):
// Xd_0__inst_mult_9_244  = SUM(( GND ) + ( Xd_0__inst_mult_9_274  ) + ( Xd_0__inst_mult_9_273  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_273 ),
	.sharein(Xd_0__inst_mult_9_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_244 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_84 (
// Equation(s):
// Xd_0__inst_mult_9_248  = SUM(( !Xd_0__inst_mult_9_272  $ (((!din_b[111]) # (!din_a[118]))) ) + ( Xd_0__inst_mult_9_278  ) + ( Xd_0__inst_mult_9_277  ))
// Xd_0__inst_mult_9_249  = CARRY(( !Xd_0__inst_mult_9_272  $ (((!din_b[111]) # (!din_a[118]))) ) + ( Xd_0__inst_mult_9_278  ) + ( Xd_0__inst_mult_9_277  ))
// Xd_0__inst_mult_9_250  = SHARE((din_b[111] & (din_a[118] & Xd_0__inst_mult_9_272 )))

	.dataa(!din_b[111]),
	.datab(!din_a[118]),
	.datac(!Xd_0__inst_mult_9_272 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_277 ),
	.sharein(Xd_0__inst_mult_9_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_248 ),
	.cout(Xd_0__inst_mult_9_249 ),
	.shareout(Xd_0__inst_mult_9_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_91 (
// Equation(s):
// Xd_0__inst_mult_14_264  = SUM(( (din_a[168] & din_b[168]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_265  = CARRY(( (din_a[168] & din_b[168]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_266  = SHARE((din_a[168] & din_b[169]))

	.dataa(!din_a[168]),
	.datab(!din_b[168]),
	.datac(!din_b[169]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_14_264 ),
	.cout(Xd_0__inst_mult_14_265 ),
	.shareout(Xd_0__inst_mult_14_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_91 (
// Equation(s):
// Xd_0__inst_mult_15_264  = SUM(( (din_a[180] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_265  = CARRY(( (din_a[180] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_266  = SHARE((din_a[180] & din_b[181]))

	.dataa(!din_a[180]),
	.datab(!din_b[180]),
	.datac(!din_b[181]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_15_264 ),
	.cout(Xd_0__inst_mult_15_265 ),
	.shareout(Xd_0__inst_mult_15_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_9 (
// Equation(s):
// Xd_0__inst_i29_9_sumout  = SUM(( !din_a[179] $ (!din_b[179]) ) + ( Xd_0__inst_mult_14_45  ) + ( Xd_0__inst_mult_14_44  ))
// Xd_0__inst_i29_10  = CARRY(( !din_a[179] $ (!din_b[179]) ) + ( Xd_0__inst_mult_14_45  ) + ( Xd_0__inst_mult_14_44  ))
// Xd_0__inst_i29_11  = SHARE(GND)

	.dataa(!din_a[179]),
	.datab(!din_b[179]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_44 ),
	.sharein(Xd_0__inst_mult_14_45 ),
	.combout(),
	.sumout(Xd_0__inst_i29_9_sumout ),
	.cout(Xd_0__inst_i29_10 ),
	.shareout(Xd_0__inst_i29_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_13 (
// Equation(s):
// Xd_0__inst_i29_13_sumout  = SUM(( !din_a[191] $ (!din_b[191]) ) + ( Xd_0__inst_i29_11  ) + ( Xd_0__inst_i29_10  ))
// Xd_0__inst_i29_14  = CARRY(( !din_a[191] $ (!din_b[191]) ) + ( Xd_0__inst_i29_11  ) + ( Xd_0__inst_i29_10  ))
// Xd_0__inst_i29_15  = SHARE(GND)

	.dataa(!din_a[191]),
	.datab(!din_b[191]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_10 ),
	.sharein(Xd_0__inst_i29_11 ),
	.combout(),
	.sumout(Xd_0__inst_i29_13_sumout ),
	.cout(Xd_0__inst_i29_14 ),
	.shareout(Xd_0__inst_i29_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_83 (
// Equation(s):
// Xd_0__inst_mult_6_244  = SUM(( GND ) + ( Xd_0__inst_mult_6_274  ) + ( Xd_0__inst_mult_6_273  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_273 ),
	.sharein(Xd_0__inst_mult_6_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_244 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_84 (
// Equation(s):
// Xd_0__inst_mult_6_248  = SUM(( !Xd_0__inst_mult_6_272  $ (((!din_b[75]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_278  ) + ( Xd_0__inst_mult_6_277  ))
// Xd_0__inst_mult_6_249  = CARRY(( !Xd_0__inst_mult_6_272  $ (((!din_b[75]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_278  ) + ( Xd_0__inst_mult_6_277  ))
// Xd_0__inst_mult_6_250  = SHARE((din_b[75] & (din_a[82] & Xd_0__inst_mult_6_272 )))

	.dataa(!din_b[75]),
	.datab(!din_a[82]),
	.datac(!Xd_0__inst_mult_6_272 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_277 ),
	.sharein(Xd_0__inst_mult_6_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_248 ),
	.cout(Xd_0__inst_mult_6_249 ),
	.shareout(Xd_0__inst_mult_6_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_92 (
// Equation(s):
// Xd_0__inst_mult_14_268  = SUM(( (!din_a[177] & (((din_a[176] & din_b[172])))) # (din_a[177] & (!din_b[171] $ (((!din_a[176]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_298  ) + ( Xd_0__inst_mult_14_297  ))
// Xd_0__inst_mult_14_269  = CARRY(( (!din_a[177] & (((din_a[176] & din_b[172])))) # (din_a[177] & (!din_b[171] $ (((!din_a[176]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_298  ) + ( Xd_0__inst_mult_14_297  ))
// Xd_0__inst_mult_14_270  = SHARE((din_a[177] & (din_b[171] & (din_a[176] & din_b[172]))))

	.dataa(!din_a[177]),
	.datab(!din_b[171]),
	.datac(!din_a[176]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_297 ),
	.sharein(Xd_0__inst_mult_14_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_268 ),
	.cout(Xd_0__inst_mult_14_269 ),
	.shareout(Xd_0__inst_mult_14_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_93 (
// Equation(s):
// Xd_0__inst_mult_14_272  = SUM(( GND ) + ( Xd_0__inst_mult_14_302  ) + ( Xd_0__inst_mult_14_301  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_301 ),
	.sharein(Xd_0__inst_mult_14_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_272 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_94 (
// Equation(s):
// Xd_0__inst_mult_14_276  = SUM(( !Xd_0__inst_mult_14_300  $ (!Xd_0__inst_mult_14_296 ) ) + ( Xd_0__inst_mult_14_306  ) + ( Xd_0__inst_mult_14_305  ))
// Xd_0__inst_mult_14_277  = CARRY(( !Xd_0__inst_mult_14_300  $ (!Xd_0__inst_mult_14_296 ) ) + ( Xd_0__inst_mult_14_306  ) + ( Xd_0__inst_mult_14_305  ))
// Xd_0__inst_mult_14_278  = SHARE((Xd_0__inst_mult_14_300  & Xd_0__inst_mult_14_296 ))

	.dataa(!Xd_0__inst_mult_14_300 ),
	.datab(!Xd_0__inst_mult_14_296 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_305 ),
	.sharein(Xd_0__inst_mult_14_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_276 ),
	.cout(Xd_0__inst_mult_14_277 ),
	.shareout(Xd_0__inst_mult_14_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_83 (
// Equation(s):
// Xd_0__inst_mult_10_244  = SUM(( (din_a[120] & din_b[120]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_245  = CARRY(( (din_a[120] & din_b[120]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_246  = SHARE((din_a[120] & din_b[121]))

	.dataa(!din_a[120]),
	.datab(!din_b[120]),
	.datac(!din_b[121]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_10_244 ),
	.cout(Xd_0__inst_mult_10_245 ),
	.shareout(Xd_0__inst_mult_10_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_87 (
// Equation(s):
// Xd_0__inst_mult_11_248  = SUM(( (din_a[132] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_249  = CARRY(( (din_a[132] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_250  = SHARE((din_a[132] & din_b[133]))

	.dataa(!din_a[132]),
	.datab(!din_b[132]),
	.datac(!din_b[133]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_248 ),
	.cout(Xd_0__inst_mult_11_249 ),
	.shareout(Xd_0__inst_mult_11_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_17 (
// Equation(s):
// Xd_0__inst_i29_17_sumout  = SUM(( !din_a[131] $ (!din_b[131]) ) + ( Xd_0__inst_i29_7  ) + ( Xd_0__inst_i29_6  ))
// Xd_0__inst_i29_18  = CARRY(( !din_a[131] $ (!din_b[131]) ) + ( Xd_0__inst_i29_7  ) + ( Xd_0__inst_i29_6  ))
// Xd_0__inst_i29_19  = SHARE(GND)

	.dataa(!din_a[131]),
	.datab(!din_b[131]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_6 ),
	.sharein(Xd_0__inst_i29_7 ),
	.combout(),
	.sumout(Xd_0__inst_i29_17_sumout ),
	.cout(Xd_0__inst_i29_18 ),
	.shareout(Xd_0__inst_i29_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_21 (
// Equation(s):
// Xd_0__inst_i29_21_sumout  = SUM(( !din_a[143] $ (!din_b[143]) ) + ( Xd_0__inst_i29_19  ) + ( Xd_0__inst_i29_18  ))
// Xd_0__inst_i29_22  = CARRY(( !din_a[143] $ (!din_b[143]) ) + ( Xd_0__inst_i29_19  ) + ( Xd_0__inst_i29_18  ))
// Xd_0__inst_i29_23  = SHARE(GND)

	.dataa(!din_a[143]),
	.datab(!din_b[143]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_18 ),
	.sharein(Xd_0__inst_i29_19 ),
	.combout(),
	.sumout(Xd_0__inst_i29_21_sumout ),
	.cout(Xd_0__inst_i29_22 ),
	.shareout(Xd_0__inst_i29_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_87 (
// Equation(s):
// Xd_0__inst_mult_8_248  = SUM(( GND ) + ( Xd_0__inst_mult_8_278  ) + ( Xd_0__inst_mult_8_277  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_277 ),
	.sharein(Xd_0__inst_mult_8_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_248 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_88 (
// Equation(s):
// Xd_0__inst_mult_8_252  = SUM(( !Xd_0__inst_mult_8_276  $ (((!din_b[99]) # (!din_a[106]))) ) + ( Xd_0__inst_mult_8_282  ) + ( Xd_0__inst_mult_8_281  ))
// Xd_0__inst_mult_8_253  = CARRY(( !Xd_0__inst_mult_8_276  $ (((!din_b[99]) # (!din_a[106]))) ) + ( Xd_0__inst_mult_8_282  ) + ( Xd_0__inst_mult_8_281  ))
// Xd_0__inst_mult_8_254  = SHARE((din_b[99] & (din_a[106] & Xd_0__inst_mult_8_276 )))

	.dataa(!din_b[99]),
	.datab(!din_a[106]),
	.datac(!Xd_0__inst_mult_8_276 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_281 ),
	.sharein(Xd_0__inst_mult_8_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_252 ),
	.cout(Xd_0__inst_mult_8_253 ),
	.shareout(Xd_0__inst_mult_8_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_89 (
// Equation(s):
// Xd_0__inst_mult_8_256  = SUM(( (din_a[96] & din_b[96]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_257  = CARRY(( (din_a[96] & din_b[96]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_258  = SHARE((din_a[96] & din_b[97]))

	.dataa(!din_a[96]),
	.datab(!din_b[96]),
	.datac(!din_b[97]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_8_256 ),
	.cout(Xd_0__inst_mult_8_257 ),
	.shareout(Xd_0__inst_mult_8_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_85 (
// Equation(s):
// Xd_0__inst_mult_9_252  = SUM(( (din_a[108] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_253  = CARRY(( (din_a[108] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_254  = SHARE((din_a[108] & din_b[109]))

	.dataa(!din_a[108]),
	.datab(!din_b[108]),
	.datac(!din_b[109]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_252 ),
	.cout(Xd_0__inst_mult_9_253 ),
	.shareout(Xd_0__inst_mult_9_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_25 (
// Equation(s):
// Xd_0__inst_i29_25_sumout  = SUM(( !din_a[107] $ (!din_b[107]) ) + ( Xd_0__inst_i29_63  ) + ( Xd_0__inst_i29_62  ))
// Xd_0__inst_i29_26  = CARRY(( !din_a[107] $ (!din_b[107]) ) + ( Xd_0__inst_i29_63  ) + ( Xd_0__inst_i29_62  ))
// Xd_0__inst_i29_27  = SHARE(GND)

	.dataa(!din_a[107]),
	.datab(!din_b[107]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_62 ),
	.sharein(Xd_0__inst_i29_63 ),
	.combout(),
	.sumout(Xd_0__inst_i29_25_sumout ),
	.cout(Xd_0__inst_i29_26 ),
	.shareout(Xd_0__inst_i29_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_29 (
// Equation(s):
// Xd_0__inst_i29_29_sumout  = SUM(( !din_a[119] $ (!din_b[119]) ) + ( Xd_0__inst_mult_9_37  ) + ( Xd_0__inst_mult_9_36  ))
// Xd_0__inst_i29_30  = CARRY(( !din_a[119] $ (!din_b[119]) ) + ( Xd_0__inst_mult_9_37  ) + ( Xd_0__inst_mult_9_36  ))
// Xd_0__inst_i29_31  = SHARE(GND)

	.dataa(!din_a[119]),
	.datab(!din_b[119]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_36 ),
	.sharein(Xd_0__inst_mult_9_37 ),
	.combout(),
	.sumout(Xd_0__inst_i29_29_sumout ),
	.cout(Xd_0__inst_i29_30 ),
	.shareout(Xd_0__inst_i29_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_88 (
// Equation(s):
// Xd_0__inst_mult_11_252  = SUM(( GND ) + ( Xd_0__inst_mult_11_278  ) + ( Xd_0__inst_mult_11_277  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_277 ),
	.sharein(Xd_0__inst_mult_11_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_252 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_89 (
// Equation(s):
// Xd_0__inst_mult_11_256  = SUM(( !Xd_0__inst_mult_11_276  $ (((!din_b[135]) # (!din_a[142]))) ) + ( Xd_0__inst_mult_11_282  ) + ( Xd_0__inst_mult_11_281  ))
// Xd_0__inst_mult_11_257  = CARRY(( !Xd_0__inst_mult_11_276  $ (((!din_b[135]) # (!din_a[142]))) ) + ( Xd_0__inst_mult_11_282  ) + ( Xd_0__inst_mult_11_281  ))
// Xd_0__inst_mult_11_258  = SHARE((din_b[135] & (din_a[142] & Xd_0__inst_mult_11_276 )))

	.dataa(!din_b[135]),
	.datab(!din_a[142]),
	.datac(!Xd_0__inst_mult_11_276 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_281 ),
	.sharein(Xd_0__inst_mult_11_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_256 ),
	.cout(Xd_0__inst_mult_11_257 ),
	.shareout(Xd_0__inst_mult_11_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_85 (
// Equation(s):
// Xd_0__inst_mult_6_252  = SUM(( (din_a[72] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_253  = CARRY(( (din_a[72] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_254  = SHARE((din_a[72] & din_b[73]))

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(!din_b[73]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_252 ),
	.cout(Xd_0__inst_mult_6_253 ),
	.shareout(Xd_0__inst_mult_6_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_81 (
// Equation(s):
// Xd_0__inst_mult_7_236  = SUM(( (din_a[84] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_237  = CARRY(( (din_a[84] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_238  = SHARE((din_a[84] & din_b[85]))

	.dataa(!din_a[84]),
	.datab(!din_b[84]),
	.datac(!din_b[85]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_236 ),
	.cout(Xd_0__inst_mult_7_237 ),
	.shareout(Xd_0__inst_mult_7_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_33 (
// Equation(s):
// Xd_0__inst_i29_33_sumout  = SUM(( !din_a[83] $ (!din_b[83]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_34  = CARRY(( !din_a[83] $ (!din_b[83]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_35  = SHARE(GND)

	.dataa(!din_a[83]),
	.datab(!din_b[83]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i29_33_sumout ),
	.cout(Xd_0__inst_i29_34 ),
	.shareout(Xd_0__inst_i29_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_37 (
// Equation(s):
// Xd_0__inst_i29_37_sumout  = SUM(( !din_a[95] $ (!din_b[95]) ) + ( Xd_0__inst_i29_35  ) + ( Xd_0__inst_i29_34  ))
// Xd_0__inst_i29_38  = CARRY(( !din_a[95] $ (!din_b[95]) ) + ( Xd_0__inst_i29_35  ) + ( Xd_0__inst_i29_34  ))
// Xd_0__inst_i29_39  = SHARE(GND)

	.dataa(!din_a[95]),
	.datab(!din_b[95]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_34 ),
	.sharein(Xd_0__inst_i29_35 ),
	.combout(),
	.sumout(Xd_0__inst_i29_37_sumout ),
	.cout(Xd_0__inst_i29_38 ),
	.shareout(Xd_0__inst_i29_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_84 (
// Equation(s):
// Xd_0__inst_mult_10_248  = SUM(( GND ) + ( Xd_0__inst_mult_10_274  ) + ( Xd_0__inst_mult_10_273  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_273 ),
	.sharein(Xd_0__inst_mult_10_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_248 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_85 (
// Equation(s):
// Xd_0__inst_mult_10_252  = SUM(( !Xd_0__inst_mult_10_272  $ (((!din_b[123]) # (!din_a[130]))) ) + ( Xd_0__inst_mult_10_278  ) + ( Xd_0__inst_mult_10_277  ))
// Xd_0__inst_mult_10_253  = CARRY(( !Xd_0__inst_mult_10_272  $ (((!din_b[123]) # (!din_a[130]))) ) + ( Xd_0__inst_mult_10_278  ) + ( Xd_0__inst_mult_10_277  ))
// Xd_0__inst_mult_10_254  = SHARE((din_b[123] & (din_a[130] & Xd_0__inst_mult_10_272 )))

	.dataa(!din_b[123]),
	.datab(!din_a[130]),
	.datac(!Xd_0__inst_mult_10_272 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_277 ),
	.sharein(Xd_0__inst_mult_10_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_252 ),
	.cout(Xd_0__inst_mult_10_253 ),
	.shareout(Xd_0__inst_mult_10_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_92 (
// Equation(s):
// Xd_0__inst_mult_15_268  = SUM(( (!din_a[187] & (((din_a[186] & din_b[189])))) # (din_a[187] & (!din_b[188] $ (((!din_a[186]) # (!din_b[189]))))) ) + ( Xd_0__inst_mult_15_298  ) + ( Xd_0__inst_mult_15_297  ))
// Xd_0__inst_mult_15_269  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[189])))) # (din_a[187] & (!din_b[188] $ (((!din_a[186]) # (!din_b[189]))))) ) + ( Xd_0__inst_mult_15_298  ) + ( Xd_0__inst_mult_15_297  ))
// Xd_0__inst_mult_15_270  = SHARE((din_a[187] & (din_b[188] & (din_a[186] & din_b[189]))))

	.dataa(!din_a[187]),
	.datab(!din_b[188]),
	.datac(!din_a[186]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_297 ),
	.sharein(Xd_0__inst_mult_15_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_268 ),
	.cout(Xd_0__inst_mult_15_269 ),
	.shareout(Xd_0__inst_mult_15_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_91 (
// Equation(s):
// Xd_0__inst_mult_4_264  = SUM(( (din_a[48] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_265  = CARRY(( (din_a[48] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_266  = SHARE((din_a[48] & din_b[49]))

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(!din_b[49]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_264 ),
	.cout(Xd_0__inst_mult_4_265 ),
	.shareout(Xd_0__inst_mult_4_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_81 (
// Equation(s):
// Xd_0__inst_mult_5_236  = SUM(( (din_a[60] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_237  = CARRY(( (din_a[60] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_238  = SHARE((din_a[60] & din_b[61]))

	.dataa(!din_a[60]),
	.datab(!din_b[60]),
	.datac(!din_b[61]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_236 ),
	.cout(Xd_0__inst_mult_5_237 ),
	.shareout(Xd_0__inst_mult_5_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_41 (
// Equation(s):
// Xd_0__inst_i29_41_sumout  = SUM(( !din_a[59] $ (!din_b[59]) ) + ( Xd_0__inst_i29_39  ) + ( Xd_0__inst_i29_38  ))
// Xd_0__inst_i29_42  = CARRY(( !din_a[59] $ (!din_b[59]) ) + ( Xd_0__inst_i29_39  ) + ( Xd_0__inst_i29_38  ))
// Xd_0__inst_i29_43  = SHARE(GND)

	.dataa(!din_a[59]),
	.datab(!din_b[59]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_38 ),
	.sharein(Xd_0__inst_i29_39 ),
	.combout(),
	.sumout(Xd_0__inst_i29_41_sumout ),
	.cout(Xd_0__inst_i29_42 ),
	.shareout(Xd_0__inst_i29_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_45 (
// Equation(s):
// Xd_0__inst_i29_45_sumout  = SUM(( !din_a[71] $ (!din_b[71]) ) + ( Xd_0__inst_i29_43  ) + ( Xd_0__inst_i29_42  ))
// Xd_0__inst_i29_46  = CARRY(( !din_a[71] $ (!din_b[71]) ) + ( Xd_0__inst_i29_43  ) + ( Xd_0__inst_i29_42  ))
// Xd_0__inst_i29_47  = SHARE(GND)

	.dataa(!din_a[71]),
	.datab(!din_b[71]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_42 ),
	.sharein(Xd_0__inst_i29_43 ),
	.combout(),
	.sumout(Xd_0__inst_i29_45_sumout ),
	.cout(Xd_0__inst_i29_46 ),
	.shareout(Xd_0__inst_i29_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_88 (
// Equation(s):
// Xd_0__inst_mult_13_252  = SUM(( GND ) + ( Xd_0__inst_mult_13_278  ) + ( Xd_0__inst_mult_13_277  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_277 ),
	.sharein(Xd_0__inst_mult_13_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_252 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_89 (
// Equation(s):
// Xd_0__inst_mult_13_256  = SUM(( !Xd_0__inst_mult_13_276  $ (((!din_b[159]) # (!din_a[166]))) ) + ( Xd_0__inst_mult_13_282  ) + ( Xd_0__inst_mult_13_281  ))
// Xd_0__inst_mult_13_257  = CARRY(( !Xd_0__inst_mult_13_276  $ (((!din_b[159]) # (!din_a[166]))) ) + ( Xd_0__inst_mult_13_282  ) + ( Xd_0__inst_mult_13_281  ))
// Xd_0__inst_mult_13_258  = SHARE((din_b[159] & (din_a[166] & Xd_0__inst_mult_13_276 )))

	.dataa(!din_b[159]),
	.datab(!din_a[166]),
	.datac(!Xd_0__inst_mult_13_276 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_281 ),
	.sharein(Xd_0__inst_mult_13_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_256 ),
	.cout(Xd_0__inst_mult_13_257 ),
	.shareout(Xd_0__inst_mult_13_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_85 (
// Equation(s):
// Xd_0__inst_mult_2_240  = SUM(( (din_a[24] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_241  = CARRY(( (din_a[24] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_242  = SHARE((din_a[24] & din_b[25]))

	.dataa(!din_a[24]),
	.datab(!din_b[24]),
	.datac(!din_b[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_240 ),
	.cout(Xd_0__inst_mult_2_241 ),
	.shareout(Xd_0__inst_mult_2_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_81 (
// Equation(s):
// Xd_0__inst_mult_3_236  = SUM(( (din_a[36] & din_b[36]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_237  = CARRY(( (din_a[36] & din_b[36]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_238  = SHARE((din_a[36] & din_b[37]))

	.dataa(!din_a[36]),
	.datab(!din_b[36]),
	.datac(!din_b[37]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_236 ),
	.cout(Xd_0__inst_mult_3_237 ),
	.shareout(Xd_0__inst_mult_3_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_49 (
// Equation(s):
// Xd_0__inst_i29_49_sumout  = SUM(( !din_a[35] $ (!din_b[35]) ) + ( Xd_0__inst_i29_47  ) + ( Xd_0__inst_i29_46  ))
// Xd_0__inst_i29_50  = CARRY(( !din_a[35] $ (!din_b[35]) ) + ( Xd_0__inst_i29_47  ) + ( Xd_0__inst_i29_46  ))
// Xd_0__inst_i29_51  = SHARE(GND)

	.dataa(!din_a[35]),
	.datab(!din_b[35]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_46 ),
	.sharein(Xd_0__inst_i29_47 ),
	.combout(),
	.sumout(Xd_0__inst_i29_49_sumout ),
	.cout(Xd_0__inst_i29_50 ),
	.shareout(Xd_0__inst_i29_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_53 (
// Equation(s):
// Xd_0__inst_i29_53_sumout  = SUM(( !din_a[47] $ (!din_b[47]) ) + ( Xd_0__inst_i29_51  ) + ( Xd_0__inst_i29_50  ))
// Xd_0__inst_i29_54  = CARRY(( !din_a[47] $ (!din_b[47]) ) + ( Xd_0__inst_i29_51  ) + ( Xd_0__inst_i29_50  ))
// Xd_0__inst_i29_55  = SHARE(GND)

	.dataa(!din_a[47]),
	.datab(!din_b[47]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_50 ),
	.sharein(Xd_0__inst_i29_51 ),
	.combout(),
	.sumout(Xd_0__inst_i29_53_sumout ),
	.cout(Xd_0__inst_i29_54 ),
	.shareout(Xd_0__inst_i29_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_93 (
// Equation(s):
// Xd_0__inst_mult_15_272  = SUM(( GND ) + ( Xd_0__inst_mult_15_302  ) + ( Xd_0__inst_mult_15_301  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_301 ),
	.sharein(Xd_0__inst_mult_15_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_272 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_94 (
// Equation(s):
// Xd_0__inst_mult_15_276  = SUM(( !Xd_0__inst_mult_15_300  $ (((!din_b[183]) # (!din_a[190]))) ) + ( Xd_0__inst_mult_15_306  ) + ( Xd_0__inst_mult_15_305  ))
// Xd_0__inst_mult_15_277  = CARRY(( !Xd_0__inst_mult_15_300  $ (((!din_b[183]) # (!din_a[190]))) ) + ( Xd_0__inst_mult_15_306  ) + ( Xd_0__inst_mult_15_305  ))
// Xd_0__inst_mult_15_278  = SHARE((din_b[183] & (din_a[190] & Xd_0__inst_mult_15_300 )))

	.dataa(!din_b[183]),
	.datab(!din_a[190]),
	.datac(!Xd_0__inst_mult_15_300 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_305 ),
	.sharein(Xd_0__inst_mult_15_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_276 ),
	.cout(Xd_0__inst_mult_15_277 ),
	.shareout(Xd_0__inst_mult_15_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_85 (
// Equation(s):
// Xd_0__inst_mult_0_240  = SUM(( (din_a[0] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_241  = CARRY(( (din_a[0] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_242  = SHARE((din_a[0] & din_b[1]))

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(!din_b[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_240 ),
	.cout(Xd_0__inst_mult_0_241 ),
	.shareout(Xd_0__inst_mult_0_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_85 (
// Equation(s):
// Xd_0__inst_mult_1_240  = SUM(( (din_a[12] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_241  = CARRY(( (din_a[12] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_242  = SHARE((din_a[12] & din_b[13]))

	.dataa(!din_a[12]),
	.datab(!din_b[12]),
	.datac(!din_b[13]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_240 ),
	.cout(Xd_0__inst_mult_1_241 ),
	.shareout(Xd_0__inst_mult_1_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_57 (
// Equation(s):
// Xd_0__inst_i29_57_sumout  = SUM(( !din_a[11] $ (!din_b[11]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_58  = CARRY(( !din_a[11] $ (!din_b[11]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_59  = SHARE(GND)

	.dataa(!din_a[11]),
	.datab(!din_b[11]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i29_57_sumout ),
	.cout(Xd_0__inst_i29_58 ),
	.shareout(Xd_0__inst_i29_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_61 (
// Equation(s):
// Xd_0__inst_i29_61_sumout  = SUM(( !din_a[23] $ (!din_b[23]) ) + ( Xd_0__inst_i29_59  ) + ( Xd_0__inst_i29_58  ))
// Xd_0__inst_i29_62  = CARRY(( !din_a[23] $ (!din_b[23]) ) + ( Xd_0__inst_i29_59  ) + ( Xd_0__inst_i29_58  ))
// Xd_0__inst_i29_63  = SHARE(GND)

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_58 ),
	.sharein(Xd_0__inst_i29_59 ),
	.combout(),
	.sumout(Xd_0__inst_i29_61_sumout ),
	.cout(Xd_0__inst_i29_62 ),
	.shareout(Xd_0__inst_i29_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_88 (
// Equation(s):
// Xd_0__inst_mult_12_264  = SUM(( GND ) + ( Xd_0__inst_mult_12_294  ) + ( Xd_0__inst_mult_12_293  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_293 ),
	.sharein(Xd_0__inst_mult_12_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_264 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_89 (
// Equation(s):
// Xd_0__inst_mult_12_268  = SUM(( !Xd_0__inst_mult_12_292  $ (((!din_b[147]) # (!din_a[154]))) ) + ( Xd_0__inst_mult_12_298  ) + ( Xd_0__inst_mult_12_297  ))
// Xd_0__inst_mult_12_269  = CARRY(( !Xd_0__inst_mult_12_292  $ (((!din_b[147]) # (!din_a[154]))) ) + ( Xd_0__inst_mult_12_298  ) + ( Xd_0__inst_mult_12_297  ))
// Xd_0__inst_mult_12_270  = SHARE((din_b[147] & (din_a[154] & Xd_0__inst_mult_12_292 )))

	.dataa(!din_b[147]),
	.datab(!din_a[154]),
	.datac(!Xd_0__inst_mult_12_292 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_297 ),
	.sharein(Xd_0__inst_mult_12_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_268 ),
	.cout(Xd_0__inst_mult_12_269 ),
	.shareout(Xd_0__inst_mult_12_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_90 (
// Equation(s):
// Xd_0__inst_mult_12_272  = SUM(( (!din_a[151] & (((din_a[150] & din_b[153])))) # (din_a[151] & (!din_b[152] $ (((!din_a[150]) # (!din_b[153]))))) ) + ( Xd_0__inst_mult_12_302  ) + ( Xd_0__inst_mult_12_301  ))
// Xd_0__inst_mult_12_273  = CARRY(( (!din_a[151] & (((din_a[150] & din_b[153])))) # (din_a[151] & (!din_b[152] $ (((!din_a[150]) # (!din_b[153]))))) ) + ( Xd_0__inst_mult_12_302  ) + ( Xd_0__inst_mult_12_301  ))
// Xd_0__inst_mult_12_274  = SHARE((din_a[151] & (din_b[152] & (din_a[150] & din_b[153]))))

	.dataa(!din_a[151]),
	.datab(!din_b[152]),
	.datac(!din_a[150]),
	.datad(!din_b[153]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_301 ),
	.sharein(Xd_0__inst_mult_12_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_272 ),
	.cout(Xd_0__inst_mult_12_273 ),
	.shareout(Xd_0__inst_mult_12_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_92 (
// Equation(s):
// Xd_0__inst_mult_4_268  = SUM(( (din_a[52] & din_b[57]) ) + ( Xd_0__inst_mult_4_290  ) + ( Xd_0__inst_mult_4_289  ))
// Xd_0__inst_mult_4_269  = CARRY(( (din_a[52] & din_b[57]) ) + ( Xd_0__inst_mult_4_290  ) + ( Xd_0__inst_mult_4_289  ))
// Xd_0__inst_mult_4_270  = SHARE((din_a[52] & din_b[58]))

	.dataa(!din_a[52]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_289 ),
	.sharein(Xd_0__inst_mult_4_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_268 ),
	.cout(Xd_0__inst_mult_4_269 ),
	.shareout(Xd_0__inst_mult_4_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_91 (
// Equation(s):
// Xd_0__inst_mult_12_276  = SUM(( (din_a[145] & din_b[144]) ) + ( Xd_0__inst_mult_12_262  ) + ( Xd_0__inst_mult_12_261  ))
// Xd_0__inst_mult_12_277  = CARRY(( (din_a[145] & din_b[144]) ) + ( Xd_0__inst_mult_12_262  ) + ( Xd_0__inst_mult_12_261  ))
// Xd_0__inst_mult_12_278  = SHARE((din_a[144] & din_b[146]))

	.dataa(!din_a[145]),
	.datab(!din_b[144]),
	.datac(!din_a[144]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_261 ),
	.sharein(Xd_0__inst_mult_12_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_276 ),
	.cout(Xd_0__inst_mult_12_277 ),
	.shareout(Xd_0__inst_mult_12_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_90 (
// Equation(s):
// Xd_0__inst_mult_13_260  = SUM(( (din_a[157] & din_b[156]) ) + ( Xd_0__inst_mult_13_250  ) + ( Xd_0__inst_mult_13_249  ))
// Xd_0__inst_mult_13_261  = CARRY(( (din_a[157] & din_b[156]) ) + ( Xd_0__inst_mult_13_250  ) + ( Xd_0__inst_mult_13_249  ))
// Xd_0__inst_mult_13_262  = SHARE((din_a[156] & din_b[158]))

	.dataa(!din_a[157]),
	.datab(!din_b[156]),
	.datac(!din_a[156]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_249 ),
	.sharein(Xd_0__inst_mult_13_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_260 ),
	.cout(Xd_0__inst_mult_13_261 ),
	.shareout(Xd_0__inst_mult_13_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_95 (
// Equation(s):
// Xd_0__inst_mult_14_280  = SUM(( (din_a[169] & din_b[168]) ) + ( Xd_0__inst_mult_14_266  ) + ( Xd_0__inst_mult_14_265  ))
// Xd_0__inst_mult_14_281  = CARRY(( (din_a[169] & din_b[168]) ) + ( Xd_0__inst_mult_14_266  ) + ( Xd_0__inst_mult_14_265  ))
// Xd_0__inst_mult_14_282  = SHARE((din_a[168] & din_b[170]))

	.dataa(!din_a[169]),
	.datab(!din_b[168]),
	.datac(!din_a[168]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_265 ),
	.sharein(Xd_0__inst_mult_14_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_280 ),
	.cout(Xd_0__inst_mult_14_281 ),
	.shareout(Xd_0__inst_mult_14_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_95 (
// Equation(s):
// Xd_0__inst_mult_15_280  = SUM(( (din_a[181] & din_b[180]) ) + ( Xd_0__inst_mult_15_266  ) + ( Xd_0__inst_mult_15_265  ))
// Xd_0__inst_mult_15_281  = CARRY(( (din_a[181] & din_b[180]) ) + ( Xd_0__inst_mult_15_266  ) + ( Xd_0__inst_mult_15_265  ))
// Xd_0__inst_mult_15_282  = SHARE((din_a[180] & din_b[182]))

	.dataa(!din_a[181]),
	.datab(!din_b[180]),
	.datac(!din_a[180]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_265 ),
	.sharein(Xd_0__inst_mult_15_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_280 ),
	.cout(Xd_0__inst_mult_15_281 ),
	.shareout(Xd_0__inst_mult_15_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_86 (
// Equation(s):
// Xd_0__inst_mult_10_256  = SUM(( (din_a[121] & din_b[120]) ) + ( Xd_0__inst_mult_10_246  ) + ( Xd_0__inst_mult_10_245  ))
// Xd_0__inst_mult_10_257  = CARRY(( (din_a[121] & din_b[120]) ) + ( Xd_0__inst_mult_10_246  ) + ( Xd_0__inst_mult_10_245  ))
// Xd_0__inst_mult_10_258  = SHARE((din_a[120] & din_b[122]))

	.dataa(!din_a[121]),
	.datab(!din_b[120]),
	.datac(!din_a[120]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_245 ),
	.sharein(Xd_0__inst_mult_10_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_256 ),
	.cout(Xd_0__inst_mult_10_257 ),
	.shareout(Xd_0__inst_mult_10_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_90 (
// Equation(s):
// Xd_0__inst_mult_11_260  = SUM(( (din_a[133] & din_b[132]) ) + ( Xd_0__inst_mult_11_250  ) + ( Xd_0__inst_mult_11_249  ))
// Xd_0__inst_mult_11_261  = CARRY(( (din_a[133] & din_b[132]) ) + ( Xd_0__inst_mult_11_250  ) + ( Xd_0__inst_mult_11_249  ))
// Xd_0__inst_mult_11_262  = SHARE((din_a[132] & din_b[134]))

	.dataa(!din_a[133]),
	.datab(!din_b[132]),
	.datac(!din_a[132]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_249 ),
	.sharein(Xd_0__inst_mult_11_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_260 ),
	.cout(Xd_0__inst_mult_11_261 ),
	.shareout(Xd_0__inst_mult_11_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_90 (
// Equation(s):
// Xd_0__inst_mult_8_260  = SUM(( (din_a[97] & din_b[96]) ) + ( Xd_0__inst_mult_8_258  ) + ( Xd_0__inst_mult_8_257  ))
// Xd_0__inst_mult_8_261  = CARRY(( (din_a[97] & din_b[96]) ) + ( Xd_0__inst_mult_8_258  ) + ( Xd_0__inst_mult_8_257  ))
// Xd_0__inst_mult_8_262  = SHARE((din_a[96] & din_b[98]))

	.dataa(!din_a[97]),
	.datab(!din_b[96]),
	.datac(!din_a[96]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_257 ),
	.sharein(Xd_0__inst_mult_8_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_260 ),
	.cout(Xd_0__inst_mult_8_261 ),
	.shareout(Xd_0__inst_mult_8_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_86 (
// Equation(s):
// Xd_0__inst_mult_9_256  = SUM(( (din_a[109] & din_b[108]) ) + ( Xd_0__inst_mult_9_254  ) + ( Xd_0__inst_mult_9_253  ))
// Xd_0__inst_mult_9_257  = CARRY(( (din_a[109] & din_b[108]) ) + ( Xd_0__inst_mult_9_254  ) + ( Xd_0__inst_mult_9_253  ))
// Xd_0__inst_mult_9_258  = SHARE((din_a[108] & din_b[110]))

	.dataa(!din_a[109]),
	.datab(!din_b[108]),
	.datac(!din_a[108]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_253 ),
	.sharein(Xd_0__inst_mult_9_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_256 ),
	.cout(Xd_0__inst_mult_9_257 ),
	.shareout(Xd_0__inst_mult_9_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_86 (
// Equation(s):
// Xd_0__inst_mult_6_256  = SUM(( (din_a[73] & din_b[72]) ) + ( Xd_0__inst_mult_6_254  ) + ( Xd_0__inst_mult_6_253  ))
// Xd_0__inst_mult_6_257  = CARRY(( (din_a[73] & din_b[72]) ) + ( Xd_0__inst_mult_6_254  ) + ( Xd_0__inst_mult_6_253  ))
// Xd_0__inst_mult_6_258  = SHARE((din_a[72] & din_b[74]))

	.dataa(!din_a[73]),
	.datab(!din_b[72]),
	.datac(!din_a[72]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_253 ),
	.sharein(Xd_0__inst_mult_6_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_256 ),
	.cout(Xd_0__inst_mult_6_257 ),
	.shareout(Xd_0__inst_mult_6_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_82 (
// Equation(s):
// Xd_0__inst_mult_7_240  = SUM(( (din_a[85] & din_b[84]) ) + ( Xd_0__inst_mult_7_238  ) + ( Xd_0__inst_mult_7_237  ))
// Xd_0__inst_mult_7_241  = CARRY(( (din_a[85] & din_b[84]) ) + ( Xd_0__inst_mult_7_238  ) + ( Xd_0__inst_mult_7_237  ))
// Xd_0__inst_mult_7_242  = SHARE((din_a[84] & din_b[86]))

	.dataa(!din_a[85]),
	.datab(!din_b[84]),
	.datac(!din_a[84]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_237 ),
	.sharein(Xd_0__inst_mult_7_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_240 ),
	.cout(Xd_0__inst_mult_7_241 ),
	.shareout(Xd_0__inst_mult_7_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_93 (
// Equation(s):
// Xd_0__inst_mult_4_272  = SUM(( (din_a[49] & din_b[48]) ) + ( Xd_0__inst_mult_4_266  ) + ( Xd_0__inst_mult_4_265  ))
// Xd_0__inst_mult_4_273  = CARRY(( (din_a[49] & din_b[48]) ) + ( Xd_0__inst_mult_4_266  ) + ( Xd_0__inst_mult_4_265  ))
// Xd_0__inst_mult_4_274  = SHARE((din_a[48] & din_b[50]))

	.dataa(!din_a[49]),
	.datab(!din_b[48]),
	.datac(!din_a[48]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_265 ),
	.sharein(Xd_0__inst_mult_4_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_272 ),
	.cout(Xd_0__inst_mult_4_273 ),
	.shareout(Xd_0__inst_mult_4_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_82 (
// Equation(s):
// Xd_0__inst_mult_5_240  = SUM(( (din_a[61] & din_b[60]) ) + ( Xd_0__inst_mult_5_238  ) + ( Xd_0__inst_mult_5_237  ))
// Xd_0__inst_mult_5_241  = CARRY(( (din_a[61] & din_b[60]) ) + ( Xd_0__inst_mult_5_238  ) + ( Xd_0__inst_mult_5_237  ))
// Xd_0__inst_mult_5_242  = SHARE((din_a[60] & din_b[62]))

	.dataa(!din_a[61]),
	.datab(!din_b[60]),
	.datac(!din_a[60]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_237 ),
	.sharein(Xd_0__inst_mult_5_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_240 ),
	.cout(Xd_0__inst_mult_5_241 ),
	.shareout(Xd_0__inst_mult_5_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_86 (
// Equation(s):
// Xd_0__inst_mult_2_244  = SUM(( (din_a[25] & din_b[24]) ) + ( Xd_0__inst_mult_2_242  ) + ( Xd_0__inst_mult_2_241  ))
// Xd_0__inst_mult_2_245  = CARRY(( (din_a[25] & din_b[24]) ) + ( Xd_0__inst_mult_2_242  ) + ( Xd_0__inst_mult_2_241  ))
// Xd_0__inst_mult_2_246  = SHARE((din_a[24] & din_b[26]))

	.dataa(!din_a[25]),
	.datab(!din_b[24]),
	.datac(!din_a[24]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_241 ),
	.sharein(Xd_0__inst_mult_2_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_244 ),
	.cout(Xd_0__inst_mult_2_245 ),
	.shareout(Xd_0__inst_mult_2_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_82 (
// Equation(s):
// Xd_0__inst_mult_3_240  = SUM(( (din_a[37] & din_b[36]) ) + ( Xd_0__inst_mult_3_238  ) + ( Xd_0__inst_mult_3_237  ))
// Xd_0__inst_mult_3_241  = CARRY(( (din_a[37] & din_b[36]) ) + ( Xd_0__inst_mult_3_238  ) + ( Xd_0__inst_mult_3_237  ))
// Xd_0__inst_mult_3_242  = SHARE((din_a[36] & din_b[38]))

	.dataa(!din_a[37]),
	.datab(!din_b[36]),
	.datac(!din_a[36]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_237 ),
	.sharein(Xd_0__inst_mult_3_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_240 ),
	.cout(Xd_0__inst_mult_3_241 ),
	.shareout(Xd_0__inst_mult_3_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_86 (
// Equation(s):
// Xd_0__inst_mult_0_244  = SUM(( (din_a[1] & din_b[0]) ) + ( Xd_0__inst_mult_0_242  ) + ( Xd_0__inst_mult_0_241  ))
// Xd_0__inst_mult_0_245  = CARRY(( (din_a[1] & din_b[0]) ) + ( Xd_0__inst_mult_0_242  ) + ( Xd_0__inst_mult_0_241  ))
// Xd_0__inst_mult_0_246  = SHARE((din_a[0] & din_b[2]))

	.dataa(!din_a[1]),
	.datab(!din_b[0]),
	.datac(!din_a[0]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_241 ),
	.sharein(Xd_0__inst_mult_0_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_244 ),
	.cout(Xd_0__inst_mult_0_245 ),
	.shareout(Xd_0__inst_mult_0_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_86 (
// Equation(s):
// Xd_0__inst_mult_1_244  = SUM(( (din_a[13] & din_b[12]) ) + ( Xd_0__inst_mult_1_242  ) + ( Xd_0__inst_mult_1_241  ))
// Xd_0__inst_mult_1_245  = CARRY(( (din_a[13] & din_b[12]) ) + ( Xd_0__inst_mult_1_242  ) + ( Xd_0__inst_mult_1_241  ))
// Xd_0__inst_mult_1_246  = SHARE((din_a[12] & din_b[14]))

	.dataa(!din_a[13]),
	.datab(!din_b[12]),
	.datac(!din_a[12]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_241 ),
	.sharein(Xd_0__inst_mult_1_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_244 ),
	.cout(Xd_0__inst_mult_1_245 ),
	.shareout(Xd_0__inst_mult_1_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_92 (
// Equation(s):
// Xd_0__inst_mult_12_280  = SUM(( (!din_a[145] & (((din_a[146] & din_b[144])))) # (din_a[145] & (!din_b[145] $ (((!din_a[146]) # (!din_b[144]))))) ) + ( Xd_0__inst_mult_12_278  ) + ( Xd_0__inst_mult_12_277  ))
// Xd_0__inst_mult_12_281  = CARRY(( (!din_a[145] & (((din_a[146] & din_b[144])))) # (din_a[145] & (!din_b[145] $ (((!din_a[146]) # (!din_b[144]))))) ) + ( Xd_0__inst_mult_12_278  ) + ( Xd_0__inst_mult_12_277  ))
// Xd_0__inst_mult_12_282  = SHARE((din_a[145] & (din_b[145] & (din_a[146] & din_b[144]))))

	.dataa(!din_a[145]),
	.datab(!din_b[145]),
	.datac(!din_a[146]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_277 ),
	.sharein(Xd_0__inst_mult_12_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_280 ),
	.cout(Xd_0__inst_mult_12_281 ),
	.shareout(Xd_0__inst_mult_12_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_91 (
// Equation(s):
// Xd_0__inst_mult_13_264  = SUM(( (!din_a[157] & (((din_a[158] & din_b[156])))) # (din_a[157] & (!din_b[157] $ (((!din_a[158]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_13_262  ) + ( Xd_0__inst_mult_13_261  ))
// Xd_0__inst_mult_13_265  = CARRY(( (!din_a[157] & (((din_a[158] & din_b[156])))) # (din_a[157] & (!din_b[157] $ (((!din_a[158]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_13_262  ) + ( Xd_0__inst_mult_13_261  ))
// Xd_0__inst_mult_13_266  = SHARE((din_a[157] & (din_b[157] & (din_a[158] & din_b[156]))))

	.dataa(!din_a[157]),
	.datab(!din_b[157]),
	.datac(!din_a[158]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_261 ),
	.sharein(Xd_0__inst_mult_13_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_264 ),
	.cout(Xd_0__inst_mult_13_265 ),
	.shareout(Xd_0__inst_mult_13_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_96 (
// Equation(s):
// Xd_0__inst_mult_14_284  = SUM(( (!din_a[169] & (((din_a[170] & din_b[168])))) # (din_a[169] & (!din_b[169] $ (((!din_a[170]) # (!din_b[168]))))) ) + ( Xd_0__inst_mult_14_282  ) + ( Xd_0__inst_mult_14_281  ))
// Xd_0__inst_mult_14_285  = CARRY(( (!din_a[169] & (((din_a[170] & din_b[168])))) # (din_a[169] & (!din_b[169] $ (((!din_a[170]) # (!din_b[168]))))) ) + ( Xd_0__inst_mult_14_282  ) + ( Xd_0__inst_mult_14_281  ))
// Xd_0__inst_mult_14_286  = SHARE((din_a[169] & (din_b[169] & (din_a[170] & din_b[168]))))

	.dataa(!din_a[169]),
	.datab(!din_b[169]),
	.datac(!din_a[170]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_281 ),
	.sharein(Xd_0__inst_mult_14_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_284 ),
	.cout(Xd_0__inst_mult_14_285 ),
	.shareout(Xd_0__inst_mult_14_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_96 (
// Equation(s):
// Xd_0__inst_mult_15_284  = SUM(( (!din_a[181] & (((din_a[182] & din_b[180])))) # (din_a[181] & (!din_b[181] $ (((!din_a[182]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_15_282  ) + ( Xd_0__inst_mult_15_281  ))
// Xd_0__inst_mult_15_285  = CARRY(( (!din_a[181] & (((din_a[182] & din_b[180])))) # (din_a[181] & (!din_b[181] $ (((!din_a[182]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_15_282  ) + ( Xd_0__inst_mult_15_281  ))
// Xd_0__inst_mult_15_286  = SHARE((din_a[181] & (din_b[181] & (din_a[182] & din_b[180]))))

	.dataa(!din_a[181]),
	.datab(!din_b[181]),
	.datac(!din_a[182]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_281 ),
	.sharein(Xd_0__inst_mult_15_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_284 ),
	.cout(Xd_0__inst_mult_15_285 ),
	.shareout(Xd_0__inst_mult_15_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_87 (
// Equation(s):
// Xd_0__inst_mult_10_260  = SUM(( (!din_a[121] & (((din_a[122] & din_b[120])))) # (din_a[121] & (!din_b[121] $ (((!din_a[122]) # (!din_b[120]))))) ) + ( Xd_0__inst_mult_10_258  ) + ( Xd_0__inst_mult_10_257  ))
// Xd_0__inst_mult_10_261  = CARRY(( (!din_a[121] & (((din_a[122] & din_b[120])))) # (din_a[121] & (!din_b[121] $ (((!din_a[122]) # (!din_b[120]))))) ) + ( Xd_0__inst_mult_10_258  ) + ( Xd_0__inst_mult_10_257  ))
// Xd_0__inst_mult_10_262  = SHARE((din_a[121] & (din_b[121] & (din_a[122] & din_b[120]))))

	.dataa(!din_a[121]),
	.datab(!din_b[121]),
	.datac(!din_a[122]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_257 ),
	.sharein(Xd_0__inst_mult_10_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_260 ),
	.cout(Xd_0__inst_mult_10_261 ),
	.shareout(Xd_0__inst_mult_10_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_91 (
// Equation(s):
// Xd_0__inst_mult_11_264  = SUM(( (!din_a[133] & (((din_a[134] & din_b[132])))) # (din_a[133] & (!din_b[133] $ (((!din_a[134]) # (!din_b[132]))))) ) + ( Xd_0__inst_mult_11_262  ) + ( Xd_0__inst_mult_11_261  ))
// Xd_0__inst_mult_11_265  = CARRY(( (!din_a[133] & (((din_a[134] & din_b[132])))) # (din_a[133] & (!din_b[133] $ (((!din_a[134]) # (!din_b[132]))))) ) + ( Xd_0__inst_mult_11_262  ) + ( Xd_0__inst_mult_11_261  ))
// Xd_0__inst_mult_11_266  = SHARE((din_a[133] & (din_b[133] & (din_a[134] & din_b[132]))))

	.dataa(!din_a[133]),
	.datab(!din_b[133]),
	.datac(!din_a[134]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_261 ),
	.sharein(Xd_0__inst_mult_11_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_264 ),
	.cout(Xd_0__inst_mult_11_265 ),
	.shareout(Xd_0__inst_mult_11_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_91 (
// Equation(s):
// Xd_0__inst_mult_8_264  = SUM(( (!din_a[97] & (((din_a[98] & din_b[96])))) # (din_a[97] & (!din_b[97] $ (((!din_a[98]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_8_262  ) + ( Xd_0__inst_mult_8_261  ))
// Xd_0__inst_mult_8_265  = CARRY(( (!din_a[97] & (((din_a[98] & din_b[96])))) # (din_a[97] & (!din_b[97] $ (((!din_a[98]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_8_262  ) + ( Xd_0__inst_mult_8_261  ))
// Xd_0__inst_mult_8_266  = SHARE((din_a[97] & (din_b[97] & (din_a[98] & din_b[96]))))

	.dataa(!din_a[97]),
	.datab(!din_b[97]),
	.datac(!din_a[98]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_261 ),
	.sharein(Xd_0__inst_mult_8_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_264 ),
	.cout(Xd_0__inst_mult_8_265 ),
	.shareout(Xd_0__inst_mult_8_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_87 (
// Equation(s):
// Xd_0__inst_mult_9_260  = SUM(( (!din_a[109] & (((din_a[110] & din_b[108])))) # (din_a[109] & (!din_b[109] $ (((!din_a[110]) # (!din_b[108]))))) ) + ( Xd_0__inst_mult_9_258  ) + ( Xd_0__inst_mult_9_257  ))
// Xd_0__inst_mult_9_261  = CARRY(( (!din_a[109] & (((din_a[110] & din_b[108])))) # (din_a[109] & (!din_b[109] $ (((!din_a[110]) # (!din_b[108]))))) ) + ( Xd_0__inst_mult_9_258  ) + ( Xd_0__inst_mult_9_257  ))
// Xd_0__inst_mult_9_262  = SHARE((din_a[109] & (din_b[109] & (din_a[110] & din_b[108]))))

	.dataa(!din_a[109]),
	.datab(!din_b[109]),
	.datac(!din_a[110]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_257 ),
	.sharein(Xd_0__inst_mult_9_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_260 ),
	.cout(Xd_0__inst_mult_9_261 ),
	.shareout(Xd_0__inst_mult_9_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_87 (
// Equation(s):
// Xd_0__inst_mult_6_260  = SUM(( (!din_a[73] & (((din_a[74] & din_b[72])))) # (din_a[73] & (!din_b[73] $ (((!din_a[74]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_258  ) + ( Xd_0__inst_mult_6_257  ))
// Xd_0__inst_mult_6_261  = CARRY(( (!din_a[73] & (((din_a[74] & din_b[72])))) # (din_a[73] & (!din_b[73] $ (((!din_a[74]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_258  ) + ( Xd_0__inst_mult_6_257  ))
// Xd_0__inst_mult_6_262  = SHARE((din_a[73] & (din_b[73] & (din_a[74] & din_b[72]))))

	.dataa(!din_a[73]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_257 ),
	.sharein(Xd_0__inst_mult_6_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_260 ),
	.cout(Xd_0__inst_mult_6_261 ),
	.shareout(Xd_0__inst_mult_6_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_83 (
// Equation(s):
// Xd_0__inst_mult_7_244  = SUM(( (!din_a[85] & (((din_a[86] & din_b[84])))) # (din_a[85] & (!din_b[85] $ (((!din_a[86]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_242  ) + ( Xd_0__inst_mult_7_241  ))
// Xd_0__inst_mult_7_245  = CARRY(( (!din_a[85] & (((din_a[86] & din_b[84])))) # (din_a[85] & (!din_b[85] $ (((!din_a[86]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_242  ) + ( Xd_0__inst_mult_7_241  ))
// Xd_0__inst_mult_7_246  = SHARE((din_a[85] & (din_b[85] & (din_a[86] & din_b[84]))))

	.dataa(!din_a[85]),
	.datab(!din_b[85]),
	.datac(!din_a[86]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_241 ),
	.sharein(Xd_0__inst_mult_7_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_244 ),
	.cout(Xd_0__inst_mult_7_245 ),
	.shareout(Xd_0__inst_mult_7_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_94 (
// Equation(s):
// Xd_0__inst_mult_4_276  = SUM(( (!din_a[49] & (((din_a[50] & din_b[48])))) # (din_a[49] & (!din_b[49] $ (((!din_a[50]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_274  ) + ( Xd_0__inst_mult_4_273  ))
// Xd_0__inst_mult_4_277  = CARRY(( (!din_a[49] & (((din_a[50] & din_b[48])))) # (din_a[49] & (!din_b[49] $ (((!din_a[50]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_274  ) + ( Xd_0__inst_mult_4_273  ))
// Xd_0__inst_mult_4_278  = SHARE((din_a[49] & (din_b[49] & (din_a[50] & din_b[48]))))

	.dataa(!din_a[49]),
	.datab(!din_b[49]),
	.datac(!din_a[50]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_273 ),
	.sharein(Xd_0__inst_mult_4_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_276 ),
	.cout(Xd_0__inst_mult_4_277 ),
	.shareout(Xd_0__inst_mult_4_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_83 (
// Equation(s):
// Xd_0__inst_mult_5_244  = SUM(( (!din_a[61] & (((din_a[62] & din_b[60])))) # (din_a[61] & (!din_b[61] $ (((!din_a[62]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_242  ) + ( Xd_0__inst_mult_5_241  ))
// Xd_0__inst_mult_5_245  = CARRY(( (!din_a[61] & (((din_a[62] & din_b[60])))) # (din_a[61] & (!din_b[61] $ (((!din_a[62]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_242  ) + ( Xd_0__inst_mult_5_241  ))
// Xd_0__inst_mult_5_246  = SHARE((din_a[61] & (din_b[61] & (din_a[62] & din_b[60]))))

	.dataa(!din_a[61]),
	.datab(!din_b[61]),
	.datac(!din_a[62]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_241 ),
	.sharein(Xd_0__inst_mult_5_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_244 ),
	.cout(Xd_0__inst_mult_5_245 ),
	.shareout(Xd_0__inst_mult_5_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_87 (
// Equation(s):
// Xd_0__inst_mult_2_248  = SUM(( (!din_a[25] & (((din_a[26] & din_b[24])))) # (din_a[25] & (!din_b[25] $ (((!din_a[26]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_246  ) + ( Xd_0__inst_mult_2_245  ))
// Xd_0__inst_mult_2_249  = CARRY(( (!din_a[25] & (((din_a[26] & din_b[24])))) # (din_a[25] & (!din_b[25] $ (((!din_a[26]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_246  ) + ( Xd_0__inst_mult_2_245  ))
// Xd_0__inst_mult_2_250  = SHARE((din_a[25] & (din_b[25] & (din_a[26] & din_b[24]))))

	.dataa(!din_a[25]),
	.datab(!din_b[25]),
	.datac(!din_a[26]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_245 ),
	.sharein(Xd_0__inst_mult_2_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_248 ),
	.cout(Xd_0__inst_mult_2_249 ),
	.shareout(Xd_0__inst_mult_2_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_83 (
// Equation(s):
// Xd_0__inst_mult_3_244  = SUM(( (!din_a[37] & (((din_a[38] & din_b[36])))) # (din_a[37] & (!din_b[37] $ (((!din_a[38]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_242  ) + ( Xd_0__inst_mult_3_241  ))
// Xd_0__inst_mult_3_245  = CARRY(( (!din_a[37] & (((din_a[38] & din_b[36])))) # (din_a[37] & (!din_b[37] $ (((!din_a[38]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_242  ) + ( Xd_0__inst_mult_3_241  ))
// Xd_0__inst_mult_3_246  = SHARE((din_a[37] & (din_b[37] & (din_a[38] & din_b[36]))))

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(!din_a[38]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_241 ),
	.sharein(Xd_0__inst_mult_3_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_244 ),
	.cout(Xd_0__inst_mult_3_245 ),
	.shareout(Xd_0__inst_mult_3_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_87 (
// Equation(s):
// Xd_0__inst_mult_0_248  = SUM(( (!din_a[1] & (((din_a[2] & din_b[0])))) # (din_a[1] & (!din_b[1] $ (((!din_a[2]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_246  ) + ( Xd_0__inst_mult_0_245  ))
// Xd_0__inst_mult_0_249  = CARRY(( (!din_a[1] & (((din_a[2] & din_b[0])))) # (din_a[1] & (!din_b[1] $ (((!din_a[2]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_246  ) + ( Xd_0__inst_mult_0_245  ))
// Xd_0__inst_mult_0_250  = SHARE((din_a[1] & (din_b[1] & (din_a[2] & din_b[0]))))

	.dataa(!din_a[1]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_245 ),
	.sharein(Xd_0__inst_mult_0_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_248 ),
	.cout(Xd_0__inst_mult_0_249 ),
	.shareout(Xd_0__inst_mult_0_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_87 (
// Equation(s):
// Xd_0__inst_mult_1_248  = SUM(( (!din_a[13] & (((din_a[14] & din_b[12])))) # (din_a[13] & (!din_b[13] $ (((!din_a[14]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_246  ) + ( Xd_0__inst_mult_1_245  ))
// Xd_0__inst_mult_1_249  = CARRY(( (!din_a[13] & (((din_a[14] & din_b[12])))) # (din_a[13] & (!din_b[13] $ (((!din_a[14]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_246  ) + ( Xd_0__inst_mult_1_245  ))
// Xd_0__inst_mult_1_250  = SHARE((din_a[13] & (din_b[13] & (din_a[14] & din_b[12]))))

	.dataa(!din_a[13]),
	.datab(!din_b[13]),
	.datac(!din_a[14]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_245 ),
	.sharein(Xd_0__inst_mult_1_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_248 ),
	.cout(Xd_0__inst_mult_1_249 ),
	.shareout(Xd_0__inst_mult_1_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_93 (
// Equation(s):
// Xd_0__inst_mult_12_284  = SUM(( (din_a[144] & din_b[147]) ) + ( Xd_0__inst_mult_12_306  ) + ( Xd_0__inst_mult_12_305  ))
// Xd_0__inst_mult_12_285  = CARRY(( (din_a[144] & din_b[147]) ) + ( Xd_0__inst_mult_12_306  ) + ( Xd_0__inst_mult_12_305  ))
// Xd_0__inst_mult_12_286  = SHARE((din_a[144] & din_b[148]))

	.dataa(!din_a[144]),
	.datab(!din_b[147]),
	.datac(!din_b[148]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_305 ),
	.sharein(Xd_0__inst_mult_12_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_284 ),
	.cout(Xd_0__inst_mult_12_285 ),
	.shareout(Xd_0__inst_mult_12_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_92 (
// Equation(s):
// Xd_0__inst_mult_13_268  = SUM(( (din_a[156] & din_b[159]) ) + ( Xd_0__inst_mult_13_286  ) + ( Xd_0__inst_mult_13_285  ))
// Xd_0__inst_mult_13_269  = CARRY(( (din_a[156] & din_b[159]) ) + ( Xd_0__inst_mult_13_286  ) + ( Xd_0__inst_mult_13_285  ))
// Xd_0__inst_mult_13_270  = SHARE((din_a[156] & din_b[160]))

	.dataa(!din_a[156]),
	.datab(!din_b[159]),
	.datac(!din_b[160]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_285 ),
	.sharein(Xd_0__inst_mult_13_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_268 ),
	.cout(Xd_0__inst_mult_13_269 ),
	.shareout(Xd_0__inst_mult_13_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_97 (
// Equation(s):
// Xd_0__inst_mult_14_288  = SUM(( (din_a[168] & din_b[171]) ) + ( Xd_0__inst_mult_14_310  ) + ( Xd_0__inst_mult_14_309  ))
// Xd_0__inst_mult_14_289  = CARRY(( (din_a[168] & din_b[171]) ) + ( Xd_0__inst_mult_14_310  ) + ( Xd_0__inst_mult_14_309  ))
// Xd_0__inst_mult_14_290  = SHARE((din_a[168] & din_b[172]))

	.dataa(!din_a[168]),
	.datab(!din_b[171]),
	.datac(!din_b[172]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_309 ),
	.sharein(Xd_0__inst_mult_14_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_288 ),
	.cout(Xd_0__inst_mult_14_289 ),
	.shareout(Xd_0__inst_mult_14_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_97 (
// Equation(s):
// Xd_0__inst_mult_15_288  = SUM(( (din_a[180] & din_b[183]) ) + ( Xd_0__inst_mult_15_310  ) + ( Xd_0__inst_mult_15_309  ))
// Xd_0__inst_mult_15_289  = CARRY(( (din_a[180] & din_b[183]) ) + ( Xd_0__inst_mult_15_310  ) + ( Xd_0__inst_mult_15_309  ))
// Xd_0__inst_mult_15_290  = SHARE((din_a[180] & din_b[184]))

	.dataa(!din_a[180]),
	.datab(!din_b[183]),
	.datac(!din_b[184]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_309 ),
	.sharein(Xd_0__inst_mult_15_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_288 ),
	.cout(Xd_0__inst_mult_15_289 ),
	.shareout(Xd_0__inst_mult_15_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_88 (
// Equation(s):
// Xd_0__inst_mult_10_264  = SUM(( (din_a[120] & din_b[123]) ) + ( Xd_0__inst_mult_10_282  ) + ( Xd_0__inst_mult_10_281  ))
// Xd_0__inst_mult_10_265  = CARRY(( (din_a[120] & din_b[123]) ) + ( Xd_0__inst_mult_10_282  ) + ( Xd_0__inst_mult_10_281  ))
// Xd_0__inst_mult_10_266  = SHARE((din_a[120] & din_b[124]))

	.dataa(!din_a[120]),
	.datab(!din_b[123]),
	.datac(!din_b[124]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_281 ),
	.sharein(Xd_0__inst_mult_10_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_264 ),
	.cout(Xd_0__inst_mult_10_265 ),
	.shareout(Xd_0__inst_mult_10_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_92 (
// Equation(s):
// Xd_0__inst_mult_11_268  = SUM(( (din_a[132] & din_b[135]) ) + ( Xd_0__inst_mult_11_286  ) + ( Xd_0__inst_mult_11_285  ))
// Xd_0__inst_mult_11_269  = CARRY(( (din_a[132] & din_b[135]) ) + ( Xd_0__inst_mult_11_286  ) + ( Xd_0__inst_mult_11_285  ))
// Xd_0__inst_mult_11_270  = SHARE((din_a[132] & din_b[136]))

	.dataa(!din_a[132]),
	.datab(!din_b[135]),
	.datac(!din_b[136]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_285 ),
	.sharein(Xd_0__inst_mult_11_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_268 ),
	.cout(Xd_0__inst_mult_11_269 ),
	.shareout(Xd_0__inst_mult_11_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_92 (
// Equation(s):
// Xd_0__inst_mult_8_268  = SUM(( (din_a[96] & din_b[99]) ) + ( Xd_0__inst_mult_8_286  ) + ( Xd_0__inst_mult_8_285  ))
// Xd_0__inst_mult_8_269  = CARRY(( (din_a[96] & din_b[99]) ) + ( Xd_0__inst_mult_8_286  ) + ( Xd_0__inst_mult_8_285  ))
// Xd_0__inst_mult_8_270  = SHARE((din_a[96] & din_b[100]))

	.dataa(!din_a[96]),
	.datab(!din_b[99]),
	.datac(!din_b[100]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_285 ),
	.sharein(Xd_0__inst_mult_8_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_268 ),
	.cout(Xd_0__inst_mult_8_269 ),
	.shareout(Xd_0__inst_mult_8_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_88 (
// Equation(s):
// Xd_0__inst_mult_9_264  = SUM(( (din_a[108] & din_b[111]) ) + ( Xd_0__inst_mult_9_282  ) + ( Xd_0__inst_mult_9_281  ))
// Xd_0__inst_mult_9_265  = CARRY(( (din_a[108] & din_b[111]) ) + ( Xd_0__inst_mult_9_282  ) + ( Xd_0__inst_mult_9_281  ))
// Xd_0__inst_mult_9_266  = SHARE((din_a[108] & din_b[112]))

	.dataa(!din_a[108]),
	.datab(!din_b[111]),
	.datac(!din_b[112]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_281 ),
	.sharein(Xd_0__inst_mult_9_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_264 ),
	.cout(Xd_0__inst_mult_9_265 ),
	.shareout(Xd_0__inst_mult_9_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_88 (
// Equation(s):
// Xd_0__inst_mult_6_264  = SUM(( (din_a[72] & din_b[75]) ) + ( Xd_0__inst_mult_6_282  ) + ( Xd_0__inst_mult_6_281  ))
// Xd_0__inst_mult_6_265  = CARRY(( (din_a[72] & din_b[75]) ) + ( Xd_0__inst_mult_6_282  ) + ( Xd_0__inst_mult_6_281  ))
// Xd_0__inst_mult_6_266  = SHARE((din_a[72] & din_b[76]))

	.dataa(!din_a[72]),
	.datab(!din_b[75]),
	.datac(!din_b[76]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_281 ),
	.sharein(Xd_0__inst_mult_6_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_264 ),
	.cout(Xd_0__inst_mult_6_265 ),
	.shareout(Xd_0__inst_mult_6_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_84 (
// Equation(s):
// Xd_0__inst_mult_7_248  = SUM(( (din_a[84] & din_b[87]) ) + ( Xd_0__inst_mult_7_258  ) + ( Xd_0__inst_mult_7_257  ))
// Xd_0__inst_mult_7_249  = CARRY(( (din_a[84] & din_b[87]) ) + ( Xd_0__inst_mult_7_258  ) + ( Xd_0__inst_mult_7_257  ))
// Xd_0__inst_mult_7_250  = SHARE((din_a[84] & din_b[88]))

	.dataa(!din_a[84]),
	.datab(!din_b[87]),
	.datac(!din_b[88]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_257 ),
	.sharein(Xd_0__inst_mult_7_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_248 ),
	.cout(Xd_0__inst_mult_7_249 ),
	.shareout(Xd_0__inst_mult_7_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_95 (
// Equation(s):
// Xd_0__inst_mult_4_280  = SUM(( (din_a[48] & din_b[51]) ) + ( Xd_0__inst_mult_4_294  ) + ( Xd_0__inst_mult_4_293  ))
// Xd_0__inst_mult_4_281  = CARRY(( (din_a[48] & din_b[51]) ) + ( Xd_0__inst_mult_4_294  ) + ( Xd_0__inst_mult_4_293  ))
// Xd_0__inst_mult_4_282  = SHARE((din_a[48] & din_b[52]))

	.dataa(!din_a[48]),
	.datab(!din_b[51]),
	.datac(!din_b[52]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_293 ),
	.sharein(Xd_0__inst_mult_4_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_280 ),
	.cout(Xd_0__inst_mult_4_281 ),
	.shareout(Xd_0__inst_mult_4_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_84 (
// Equation(s):
// Xd_0__inst_mult_5_248  = SUM(( (din_a[60] & din_b[63]) ) + ( Xd_0__inst_mult_5_258  ) + ( Xd_0__inst_mult_5_257  ))
// Xd_0__inst_mult_5_249  = CARRY(( (din_a[60] & din_b[63]) ) + ( Xd_0__inst_mult_5_258  ) + ( Xd_0__inst_mult_5_257  ))
// Xd_0__inst_mult_5_250  = SHARE((din_a[60] & din_b[64]))

	.dataa(!din_a[60]),
	.datab(!din_b[63]),
	.datac(!din_b[64]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_257 ),
	.sharein(Xd_0__inst_mult_5_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_248 ),
	.cout(Xd_0__inst_mult_5_249 ),
	.shareout(Xd_0__inst_mult_5_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_88 (
// Equation(s):
// Xd_0__inst_mult_2_252  = SUM(( (din_a[24] & din_b[27]) ) + ( Xd_0__inst_mult_2_262  ) + ( Xd_0__inst_mult_2_261  ))
// Xd_0__inst_mult_2_253  = CARRY(( (din_a[24] & din_b[27]) ) + ( Xd_0__inst_mult_2_262  ) + ( Xd_0__inst_mult_2_261  ))
// Xd_0__inst_mult_2_254  = SHARE((din_a[24] & din_b[28]))

	.dataa(!din_a[24]),
	.datab(!din_b[27]),
	.datac(!din_b[28]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_261 ),
	.sharein(Xd_0__inst_mult_2_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_252 ),
	.cout(Xd_0__inst_mult_2_253 ),
	.shareout(Xd_0__inst_mult_2_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_84 (
// Equation(s):
// Xd_0__inst_mult_3_248  = SUM(( (din_a[36] & din_b[39]) ) + ( Xd_0__inst_mult_3_258  ) + ( Xd_0__inst_mult_3_257  ))
// Xd_0__inst_mult_3_249  = CARRY(( (din_a[36] & din_b[39]) ) + ( Xd_0__inst_mult_3_258  ) + ( Xd_0__inst_mult_3_257  ))
// Xd_0__inst_mult_3_250  = SHARE((din_a[36] & din_b[40]))

	.dataa(!din_a[36]),
	.datab(!din_b[39]),
	.datac(!din_b[40]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_257 ),
	.sharein(Xd_0__inst_mult_3_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_248 ),
	.cout(Xd_0__inst_mult_3_249 ),
	.shareout(Xd_0__inst_mult_3_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_88 (
// Equation(s):
// Xd_0__inst_mult_0_252  = SUM(( (din_a[0] & din_b[3]) ) + ( Xd_0__inst_mult_0_262  ) + ( Xd_0__inst_mult_0_261  ))
// Xd_0__inst_mult_0_253  = CARRY(( (din_a[0] & din_b[3]) ) + ( Xd_0__inst_mult_0_262  ) + ( Xd_0__inst_mult_0_261  ))
// Xd_0__inst_mult_0_254  = SHARE((din_a[0] & din_b[4]))

	.dataa(!din_a[0]),
	.datab(!din_b[3]),
	.datac(!din_b[4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_261 ),
	.sharein(Xd_0__inst_mult_0_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_252 ),
	.cout(Xd_0__inst_mult_0_253 ),
	.shareout(Xd_0__inst_mult_0_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_88 (
// Equation(s):
// Xd_0__inst_mult_1_252  = SUM(( (din_a[12] & din_b[15]) ) + ( Xd_0__inst_mult_1_262  ) + ( Xd_0__inst_mult_1_261  ))
// Xd_0__inst_mult_1_253  = CARRY(( (din_a[12] & din_b[15]) ) + ( Xd_0__inst_mult_1_262  ) + ( Xd_0__inst_mult_1_261  ))
// Xd_0__inst_mult_1_254  = SHARE((din_a[12] & din_b[16]))

	.dataa(!din_a[12]),
	.datab(!din_b[15]),
	.datac(!din_b[16]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_261 ),
	.sharein(Xd_0__inst_mult_1_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_252 ),
	.cout(Xd_0__inst_mult_1_253 ),
	.shareout(Xd_0__inst_mult_1_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_94 (
// Equation(s):
// Xd_0__inst_mult_12_288  = SUM(( !Xd_0__inst_mult_12_308  $ (!Xd_0__inst_mult_12_312 ) ) + ( Xd_0__inst_mult_12_286  ) + ( Xd_0__inst_mult_12_285  ))
// Xd_0__inst_mult_12_289  = CARRY(( !Xd_0__inst_mult_12_308  $ (!Xd_0__inst_mult_12_312 ) ) + ( Xd_0__inst_mult_12_286  ) + ( Xd_0__inst_mult_12_285  ))
// Xd_0__inst_mult_12_290  = SHARE((Xd_0__inst_mult_12_308  & Xd_0__inst_mult_12_312 ))

	.dataa(!Xd_0__inst_mult_12_308 ),
	.datab(!Xd_0__inst_mult_12_312 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_285 ),
	.sharein(Xd_0__inst_mult_12_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_288 ),
	.cout(Xd_0__inst_mult_12_289 ),
	.shareout(Xd_0__inst_mult_12_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_93 (
// Equation(s):
// Xd_0__inst_mult_13_272  = SUM(( !Xd_0__inst_mult_13_288  $ (!Xd_0__inst_mult_13_292 ) ) + ( Xd_0__inst_mult_13_270  ) + ( Xd_0__inst_mult_13_269  ))
// Xd_0__inst_mult_13_273  = CARRY(( !Xd_0__inst_mult_13_288  $ (!Xd_0__inst_mult_13_292 ) ) + ( Xd_0__inst_mult_13_270  ) + ( Xd_0__inst_mult_13_269  ))
// Xd_0__inst_mult_13_274  = SHARE((Xd_0__inst_mult_13_288  & Xd_0__inst_mult_13_292 ))

	.dataa(!Xd_0__inst_mult_13_288 ),
	.datab(!Xd_0__inst_mult_13_292 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_269 ),
	.sharein(Xd_0__inst_mult_13_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_272 ),
	.cout(Xd_0__inst_mult_13_273 ),
	.shareout(Xd_0__inst_mult_13_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_98 (
// Equation(s):
// Xd_0__inst_mult_14_292  = SUM(( !Xd_0__inst_mult_14_312  $ (!Xd_0__inst_mult_14_316 ) ) + ( Xd_0__inst_mult_14_290  ) + ( Xd_0__inst_mult_14_289  ))
// Xd_0__inst_mult_14_293  = CARRY(( !Xd_0__inst_mult_14_312  $ (!Xd_0__inst_mult_14_316 ) ) + ( Xd_0__inst_mult_14_290  ) + ( Xd_0__inst_mult_14_289  ))
// Xd_0__inst_mult_14_294  = SHARE((Xd_0__inst_mult_14_312  & Xd_0__inst_mult_14_316 ))

	.dataa(!Xd_0__inst_mult_14_312 ),
	.datab(!Xd_0__inst_mult_14_316 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_289 ),
	.sharein(Xd_0__inst_mult_14_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_292 ),
	.cout(Xd_0__inst_mult_14_293 ),
	.shareout(Xd_0__inst_mult_14_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_98 (
// Equation(s):
// Xd_0__inst_mult_15_292  = SUM(( !Xd_0__inst_mult_15_312  $ (!Xd_0__inst_mult_15_316 ) ) + ( Xd_0__inst_mult_15_290  ) + ( Xd_0__inst_mult_15_289  ))
// Xd_0__inst_mult_15_293  = CARRY(( !Xd_0__inst_mult_15_312  $ (!Xd_0__inst_mult_15_316 ) ) + ( Xd_0__inst_mult_15_290  ) + ( Xd_0__inst_mult_15_289  ))
// Xd_0__inst_mult_15_294  = SHARE((Xd_0__inst_mult_15_312  & Xd_0__inst_mult_15_316 ))

	.dataa(!Xd_0__inst_mult_15_312 ),
	.datab(!Xd_0__inst_mult_15_316 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_289 ),
	.sharein(Xd_0__inst_mult_15_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_292 ),
	.cout(Xd_0__inst_mult_15_293 ),
	.shareout(Xd_0__inst_mult_15_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_89 (
// Equation(s):
// Xd_0__inst_mult_10_268  = SUM(( !Xd_0__inst_mult_10_284  $ (!Xd_0__inst_mult_10_288 ) ) + ( Xd_0__inst_mult_10_266  ) + ( Xd_0__inst_mult_10_265  ))
// Xd_0__inst_mult_10_269  = CARRY(( !Xd_0__inst_mult_10_284  $ (!Xd_0__inst_mult_10_288 ) ) + ( Xd_0__inst_mult_10_266  ) + ( Xd_0__inst_mult_10_265  ))
// Xd_0__inst_mult_10_270  = SHARE((Xd_0__inst_mult_10_284  & Xd_0__inst_mult_10_288 ))

	.dataa(!Xd_0__inst_mult_10_284 ),
	.datab(!Xd_0__inst_mult_10_288 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_265 ),
	.sharein(Xd_0__inst_mult_10_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_268 ),
	.cout(Xd_0__inst_mult_10_269 ),
	.shareout(Xd_0__inst_mult_10_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_93 (
// Equation(s):
// Xd_0__inst_mult_11_272  = SUM(( !Xd_0__inst_mult_11_288  $ (!Xd_0__inst_mult_11_292 ) ) + ( Xd_0__inst_mult_11_270  ) + ( Xd_0__inst_mult_11_269  ))
// Xd_0__inst_mult_11_273  = CARRY(( !Xd_0__inst_mult_11_288  $ (!Xd_0__inst_mult_11_292 ) ) + ( Xd_0__inst_mult_11_270  ) + ( Xd_0__inst_mult_11_269  ))
// Xd_0__inst_mult_11_274  = SHARE((Xd_0__inst_mult_11_288  & Xd_0__inst_mult_11_292 ))

	.dataa(!Xd_0__inst_mult_11_288 ),
	.datab(!Xd_0__inst_mult_11_292 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_269 ),
	.sharein(Xd_0__inst_mult_11_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_272 ),
	.cout(Xd_0__inst_mult_11_273 ),
	.shareout(Xd_0__inst_mult_11_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_93 (
// Equation(s):
// Xd_0__inst_mult_8_272  = SUM(( !Xd_0__inst_mult_8_288  $ (!Xd_0__inst_mult_8_292 ) ) + ( Xd_0__inst_mult_8_270  ) + ( Xd_0__inst_mult_8_269  ))
// Xd_0__inst_mult_8_273  = CARRY(( !Xd_0__inst_mult_8_288  $ (!Xd_0__inst_mult_8_292 ) ) + ( Xd_0__inst_mult_8_270  ) + ( Xd_0__inst_mult_8_269  ))
// Xd_0__inst_mult_8_274  = SHARE((Xd_0__inst_mult_8_288  & Xd_0__inst_mult_8_292 ))

	.dataa(!Xd_0__inst_mult_8_288 ),
	.datab(!Xd_0__inst_mult_8_292 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_269 ),
	.sharein(Xd_0__inst_mult_8_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_272 ),
	.cout(Xd_0__inst_mult_8_273 ),
	.shareout(Xd_0__inst_mult_8_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_89 (
// Equation(s):
// Xd_0__inst_mult_9_268  = SUM(( !Xd_0__inst_mult_9_284  $ (!Xd_0__inst_mult_9_288 ) ) + ( Xd_0__inst_mult_9_266  ) + ( Xd_0__inst_mult_9_265  ))
// Xd_0__inst_mult_9_269  = CARRY(( !Xd_0__inst_mult_9_284  $ (!Xd_0__inst_mult_9_288 ) ) + ( Xd_0__inst_mult_9_266  ) + ( Xd_0__inst_mult_9_265  ))
// Xd_0__inst_mult_9_270  = SHARE((Xd_0__inst_mult_9_284  & Xd_0__inst_mult_9_288 ))

	.dataa(!Xd_0__inst_mult_9_284 ),
	.datab(!Xd_0__inst_mult_9_288 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_265 ),
	.sharein(Xd_0__inst_mult_9_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_268 ),
	.cout(Xd_0__inst_mult_9_269 ),
	.shareout(Xd_0__inst_mult_9_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_89 (
// Equation(s):
// Xd_0__inst_mult_6_268  = SUM(( !Xd_0__inst_mult_6_284  $ (!Xd_0__inst_mult_6_288 ) ) + ( Xd_0__inst_mult_6_266  ) + ( Xd_0__inst_mult_6_265  ))
// Xd_0__inst_mult_6_269  = CARRY(( !Xd_0__inst_mult_6_284  $ (!Xd_0__inst_mult_6_288 ) ) + ( Xd_0__inst_mult_6_266  ) + ( Xd_0__inst_mult_6_265  ))
// Xd_0__inst_mult_6_270  = SHARE((Xd_0__inst_mult_6_284  & Xd_0__inst_mult_6_288 ))

	.dataa(!Xd_0__inst_mult_6_284 ),
	.datab(!Xd_0__inst_mult_6_288 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_265 ),
	.sharein(Xd_0__inst_mult_6_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_268 ),
	.cout(Xd_0__inst_mult_6_269 ),
	.shareout(Xd_0__inst_mult_6_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_85 (
// Equation(s):
// Xd_0__inst_mult_7_252  = SUM(( !Xd_0__inst_mult_7_260  $ (!Xd_0__inst_mult_7_264 ) ) + ( Xd_0__inst_mult_7_250  ) + ( Xd_0__inst_mult_7_249  ))
// Xd_0__inst_mult_7_253  = CARRY(( !Xd_0__inst_mult_7_260  $ (!Xd_0__inst_mult_7_264 ) ) + ( Xd_0__inst_mult_7_250  ) + ( Xd_0__inst_mult_7_249  ))
// Xd_0__inst_mult_7_254  = SHARE((Xd_0__inst_mult_7_260  & Xd_0__inst_mult_7_264 ))

	.dataa(!Xd_0__inst_mult_7_260 ),
	.datab(!Xd_0__inst_mult_7_264 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_249 ),
	.sharein(Xd_0__inst_mult_7_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_252 ),
	.cout(Xd_0__inst_mult_7_253 ),
	.shareout(Xd_0__inst_mult_7_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_96 (
// Equation(s):
// Xd_0__inst_mult_4_284  = SUM(( !Xd_0__inst_mult_4_296  $ (!Xd_0__inst_mult_4_300 ) ) + ( Xd_0__inst_mult_4_282  ) + ( Xd_0__inst_mult_4_281  ))
// Xd_0__inst_mult_4_285  = CARRY(( !Xd_0__inst_mult_4_296  $ (!Xd_0__inst_mult_4_300 ) ) + ( Xd_0__inst_mult_4_282  ) + ( Xd_0__inst_mult_4_281  ))
// Xd_0__inst_mult_4_286  = SHARE((Xd_0__inst_mult_4_296  & Xd_0__inst_mult_4_300 ))

	.dataa(!Xd_0__inst_mult_4_296 ),
	.datab(!Xd_0__inst_mult_4_300 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_281 ),
	.sharein(Xd_0__inst_mult_4_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_284 ),
	.cout(Xd_0__inst_mult_4_285 ),
	.shareout(Xd_0__inst_mult_4_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_85 (
// Equation(s):
// Xd_0__inst_mult_5_252  = SUM(( !Xd_0__inst_mult_5_260  $ (!Xd_0__inst_mult_5_264 ) ) + ( Xd_0__inst_mult_5_250  ) + ( Xd_0__inst_mult_5_249  ))
// Xd_0__inst_mult_5_253  = CARRY(( !Xd_0__inst_mult_5_260  $ (!Xd_0__inst_mult_5_264 ) ) + ( Xd_0__inst_mult_5_250  ) + ( Xd_0__inst_mult_5_249  ))
// Xd_0__inst_mult_5_254  = SHARE((Xd_0__inst_mult_5_260  & Xd_0__inst_mult_5_264 ))

	.dataa(!Xd_0__inst_mult_5_260 ),
	.datab(!Xd_0__inst_mult_5_264 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_249 ),
	.sharein(Xd_0__inst_mult_5_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_252 ),
	.cout(Xd_0__inst_mult_5_253 ),
	.shareout(Xd_0__inst_mult_5_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_89 (
// Equation(s):
// Xd_0__inst_mult_2_256  = SUM(( !Xd_0__inst_mult_2_264  $ (!Xd_0__inst_mult_2_268 ) ) + ( Xd_0__inst_mult_2_254  ) + ( Xd_0__inst_mult_2_253  ))
// Xd_0__inst_mult_2_257  = CARRY(( !Xd_0__inst_mult_2_264  $ (!Xd_0__inst_mult_2_268 ) ) + ( Xd_0__inst_mult_2_254  ) + ( Xd_0__inst_mult_2_253  ))
// Xd_0__inst_mult_2_258  = SHARE((Xd_0__inst_mult_2_264  & Xd_0__inst_mult_2_268 ))

	.dataa(!Xd_0__inst_mult_2_264 ),
	.datab(!Xd_0__inst_mult_2_268 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_253 ),
	.sharein(Xd_0__inst_mult_2_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_256 ),
	.cout(Xd_0__inst_mult_2_257 ),
	.shareout(Xd_0__inst_mult_2_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_85 (
// Equation(s):
// Xd_0__inst_mult_3_252  = SUM(( !Xd_0__inst_mult_3_260  $ (!Xd_0__inst_mult_3_264 ) ) + ( Xd_0__inst_mult_3_250  ) + ( Xd_0__inst_mult_3_249  ))
// Xd_0__inst_mult_3_253  = CARRY(( !Xd_0__inst_mult_3_260  $ (!Xd_0__inst_mult_3_264 ) ) + ( Xd_0__inst_mult_3_250  ) + ( Xd_0__inst_mult_3_249  ))
// Xd_0__inst_mult_3_254  = SHARE((Xd_0__inst_mult_3_260  & Xd_0__inst_mult_3_264 ))

	.dataa(!Xd_0__inst_mult_3_260 ),
	.datab(!Xd_0__inst_mult_3_264 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_249 ),
	.sharein(Xd_0__inst_mult_3_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_252 ),
	.cout(Xd_0__inst_mult_3_253 ),
	.shareout(Xd_0__inst_mult_3_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_89 (
// Equation(s):
// Xd_0__inst_mult_0_256  = SUM(( !Xd_0__inst_mult_0_264  $ (!Xd_0__inst_mult_0_268 ) ) + ( Xd_0__inst_mult_0_254  ) + ( Xd_0__inst_mult_0_253  ))
// Xd_0__inst_mult_0_257  = CARRY(( !Xd_0__inst_mult_0_264  $ (!Xd_0__inst_mult_0_268 ) ) + ( Xd_0__inst_mult_0_254  ) + ( Xd_0__inst_mult_0_253  ))
// Xd_0__inst_mult_0_258  = SHARE((Xd_0__inst_mult_0_264  & Xd_0__inst_mult_0_268 ))

	.dataa(!Xd_0__inst_mult_0_264 ),
	.datab(!Xd_0__inst_mult_0_268 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_253 ),
	.sharein(Xd_0__inst_mult_0_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_256 ),
	.cout(Xd_0__inst_mult_0_257 ),
	.shareout(Xd_0__inst_mult_0_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_89 (
// Equation(s):
// Xd_0__inst_mult_1_256  = SUM(( !Xd_0__inst_mult_1_264  $ (!Xd_0__inst_mult_1_268 ) ) + ( Xd_0__inst_mult_1_254  ) + ( Xd_0__inst_mult_1_253  ))
// Xd_0__inst_mult_1_257  = CARRY(( !Xd_0__inst_mult_1_264  $ (!Xd_0__inst_mult_1_268 ) ) + ( Xd_0__inst_mult_1_254  ) + ( Xd_0__inst_mult_1_253  ))
// Xd_0__inst_mult_1_258  = SHARE((Xd_0__inst_mult_1_264  & Xd_0__inst_mult_1_268 ))

	.dataa(!Xd_0__inst_mult_1_264 ),
	.datab(!Xd_0__inst_mult_1_268 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_253 ),
	.sharein(Xd_0__inst_mult_1_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_256 ),
	.cout(Xd_0__inst_mult_1_257 ),
	.shareout(Xd_0__inst_mult_1_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_35 (
// Equation(s):
// Xd_0__inst_mult_12_35_sumout  = SUM(( (din_a[154] & din_b[144]) ) + ( Xd_0__inst_mult_13_41  ) + ( Xd_0__inst_mult_13_40  ))
// Xd_0__inst_mult_12_36  = CARRY(( (din_a[154] & din_b[144]) ) + ( Xd_0__inst_mult_13_41  ) + ( Xd_0__inst_mult_13_40  ))
// Xd_0__inst_mult_12_37  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[144]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_40 ),
	.sharein(Xd_0__inst_mult_13_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_35_sumout ),
	.cout(Xd_0__inst_mult_12_36 ),
	.shareout(Xd_0__inst_mult_12_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_35 (
// Equation(s):
// Xd_0__inst_mult_1_35_sumout  = SUM(( (din_a[21] & din_b[12]) ) + ( Xd_0__inst_mult_14_49  ) + ( Xd_0__inst_mult_14_48  ))
// Xd_0__inst_mult_1_36  = CARRY(( (din_a[21] & din_b[12]) ) + ( Xd_0__inst_mult_14_49  ) + ( Xd_0__inst_mult_14_48  ))
// Xd_0__inst_mult_1_37  = SHARE(GND)

	.dataa(!din_a[21]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_48 ),
	.sharein(Xd_0__inst_mult_14_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_35_sumout ),
	.cout(Xd_0__inst_mult_1_36 ),
	.shareout(Xd_0__inst_mult_1_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_35 (
// Equation(s):
// Xd_0__inst_mult_6_35_sumout  = SUM(( (din_a[82] & din_b[72]) ) + ( Xd_0__inst_mult_7_37  ) + ( Xd_0__inst_mult_7_36  ))
// Xd_0__inst_mult_6_36  = CARRY(( (din_a[82] & din_b[72]) ) + ( Xd_0__inst_mult_7_37  ) + ( Xd_0__inst_mult_7_36  ))
// Xd_0__inst_mult_6_37  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_36 ),
	.sharein(Xd_0__inst_mult_7_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_35_sumout ),
	.cout(Xd_0__inst_mult_6_36 ),
	.shareout(Xd_0__inst_mult_6_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_35 (
// Equation(s):
// Xd_0__inst_mult_5_35_sumout  = SUM(( (din_a[69] & din_b[60]) ) + ( Xd_0__inst_mult_8_37  ) + ( Xd_0__inst_mult_8_36  ))
// Xd_0__inst_mult_5_36  = CARRY(( (din_a[69] & din_b[60]) ) + ( Xd_0__inst_mult_8_37  ) + ( Xd_0__inst_mult_8_36  ))
// Xd_0__inst_mult_5_37  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_36 ),
	.sharein(Xd_0__inst_mult_8_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_35_sumout ),
	.cout(Xd_0__inst_mult_5_36 ),
	.shareout(Xd_0__inst_mult_5_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_35 (
// Equation(s):
// Xd_0__inst_mult_2_35_sumout  = SUM(( (din_a[33] & din_b[24]) ) + ( Xd_0__inst_mult_3_41  ) + ( Xd_0__inst_mult_3_40  ))
// Xd_0__inst_mult_2_36  = CARRY(( (din_a[33] & din_b[24]) ) + ( Xd_0__inst_mult_3_41  ) + ( Xd_0__inst_mult_3_40  ))
// Xd_0__inst_mult_2_37  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_40 ),
	.sharein(Xd_0__inst_mult_3_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_35_sumout ),
	.cout(Xd_0__inst_mult_2_36 ),
	.shareout(Xd_0__inst_mult_2_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_35 (
// Equation(s):
// Xd_0__inst_mult_14_35_sumout  = SUM(( (din_a[175] & din_b[168]) ) + ( Xd_0__inst_mult_15_41  ) + ( Xd_0__inst_mult_15_40  ))
// Xd_0__inst_mult_14_36  = CARRY(( (din_a[175] & din_b[168]) ) + ( Xd_0__inst_mult_15_41  ) + ( Xd_0__inst_mult_15_40  ))
// Xd_0__inst_mult_14_37  = SHARE(GND)

	.dataa(!din_a[175]),
	.datab(!din_b[168]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_40 ),
	.sharein(Xd_0__inst_mult_15_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_35_sumout ),
	.cout(Xd_0__inst_mult_14_36 ),
	.shareout(Xd_0__inst_mult_14_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_39 (
// Equation(s):
// Xd_0__inst_mult_12_39_sumout  = SUM(( (din_a[154] & din_b[154]) ) + ( Xd_0__inst_mult_3_45  ) + ( Xd_0__inst_mult_3_44  ))
// Xd_0__inst_mult_12_40  = CARRY(( (din_a[154] & din_b[154]) ) + ( Xd_0__inst_mult_3_45  ) + ( Xd_0__inst_mult_3_44  ))
// Xd_0__inst_mult_12_41  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[154]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_44 ),
	.sharein(Xd_0__inst_mult_3_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_39_sumout ),
	.cout(Xd_0__inst_mult_12_40 ),
	.shareout(Xd_0__inst_mult_12_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_35 (
// Equation(s):
// Xd_0__inst_mult_15_35_sumout  = SUM(( (din_a[190] & din_b[190]) ) + ( Xd_0__inst_mult_1_41  ) + ( Xd_0__inst_mult_1_40  ))
// Xd_0__inst_mult_15_36  = CARRY(( (din_a[190] & din_b[190]) ) + ( Xd_0__inst_mult_1_41  ) + ( Xd_0__inst_mult_1_40  ))
// Xd_0__inst_mult_15_37  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[190]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_40 ),
	.sharein(Xd_0__inst_mult_1_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_35_sumout ),
	.cout(Xd_0__inst_mult_15_36 ),
	.shareout(Xd_0__inst_mult_15_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_39 (
// Equation(s):
// Xd_0__inst_mult_5_39_sumout  = SUM(( (din_a[70] & din_b[70]) ) + ( Xd_0__inst_mult_12_45  ) + ( Xd_0__inst_mult_12_44  ))
// Xd_0__inst_mult_5_40  = CARRY(( (din_a[70] & din_b[70]) ) + ( Xd_0__inst_mult_12_45  ) + ( Xd_0__inst_mult_12_44  ))
// Xd_0__inst_mult_5_41  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_44 ),
	.sharein(Xd_0__inst_mult_12_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_39_sumout ),
	.cout(Xd_0__inst_mult_5_40 ),
	.shareout(Xd_0__inst_mult_5_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_35 (
// Equation(s):
// Xd_0__inst_mult_4_35_sumout  = SUM(( (din_a[58] & din_b[58]) ) + ( Xd_0__inst_mult_11_37  ) + ( Xd_0__inst_mult_11_36  ))
// Xd_0__inst_mult_4_36  = CARRY(( (din_a[58] & din_b[58]) ) + ( Xd_0__inst_mult_11_37  ) + ( Xd_0__inst_mult_11_36  ))
// Xd_0__inst_mult_4_37  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_36 ),
	.sharein(Xd_0__inst_mult_11_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_35_sumout ),
	.cout(Xd_0__inst_mult_4_36 ),
	.shareout(Xd_0__inst_mult_4_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_35 (
// Equation(s):
// Xd_0__inst_mult_10_35_sumout  = SUM(( (din_a[127] & din_b[120]) ) + ( Xd_0__inst_mult_8_41  ) + ( Xd_0__inst_mult_8_40  ))
// Xd_0__inst_mult_10_36  = CARRY(( (din_a[127] & din_b[120]) ) + ( Xd_0__inst_mult_8_41  ) + ( Xd_0__inst_mult_8_40  ))
// Xd_0__inst_mult_10_37  = SHARE(GND)

	.dataa(!din_a[127]),
	.datab(!din_b[120]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_40 ),
	.sharein(Xd_0__inst_mult_8_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_35_sumout ),
	.cout(Xd_0__inst_mult_10_36 ),
	.shareout(Xd_0__inst_mult_10_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_39 (
// Equation(s):
// Xd_0__inst_mult_6_39_sumout  = SUM(( (din_a[82] & din_b[82]) ) + ( Xd_0__inst_mult_8_45  ) + ( Xd_0__inst_mult_8_44  ))
// Xd_0__inst_mult_6_40  = CARRY(( (din_a[82] & din_b[82]) ) + ( Xd_0__inst_mult_8_45  ) + ( Xd_0__inst_mult_8_44  ))
// Xd_0__inst_mult_6_41  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_44 ),
	.sharein(Xd_0__inst_mult_8_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_39_sumout ),
	.cout(Xd_0__inst_mult_6_40 ),
	.shareout(Xd_0__inst_mult_6_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_39 (
// Equation(s):
// Xd_0__inst_mult_2_39_sumout  = SUM(( (din_a[34] & din_b[34]) ) + ( Xd_0__inst_mult_14_53  ) + ( Xd_0__inst_mult_14_52  ))
// Xd_0__inst_mult_2_40  = CARRY(( (din_a[34] & din_b[34]) ) + ( Xd_0__inst_mult_14_53  ) + ( Xd_0__inst_mult_14_52  ))
// Xd_0__inst_mult_2_41  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_52 ),
	.sharein(Xd_0__inst_mult_14_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_39_sumout ),
	.cout(Xd_0__inst_mult_2_40 ),
	.shareout(Xd_0__inst_mult_2_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_35 (
// Equation(s):
// Xd_0__inst_mult_13_35_sumout  = SUM(( (din_a[164] & din_b[156]) ) + ( Xd_0__inst_mult_10_41  ) + ( Xd_0__inst_mult_10_40  ))
// Xd_0__inst_mult_13_36  = CARRY(( (din_a[164] & din_b[156]) ) + ( Xd_0__inst_mult_10_41  ) + ( Xd_0__inst_mult_10_40  ))
// Xd_0__inst_mult_13_37  = SHARE(GND)

	.dataa(!din_a[164]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_40 ),
	.sharein(Xd_0__inst_mult_10_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_35_sumout ),
	.cout(Xd_0__inst_mult_13_36 ),
	.shareout(Xd_0__inst_mult_13_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_39 (
// Equation(s):
// Xd_0__inst_mult_14_39_sumout  = SUM(( (din_a[176] & din_b[168]) ) + ( Xd_0__inst_mult_15_45  ) + ( Xd_0__inst_mult_15_44  ))
// Xd_0__inst_mult_14_40  = CARRY(( (din_a[176] & din_b[168]) ) + ( Xd_0__inst_mult_15_45  ) + ( Xd_0__inst_mult_15_44  ))
// Xd_0__inst_mult_14_41  = SHARE(GND)

	.dataa(!din_a[176]),
	.datab(!din_b[168]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_44 ),
	.sharein(Xd_0__inst_mult_15_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_39_sumout ),
	.cout(Xd_0__inst_mult_14_40 ),
	.shareout(Xd_0__inst_mult_14_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_35 (
// Equation(s):
// Xd_0__inst_mult_3_35_sumout  = SUM(( (din_a[43] & din_b[36]) ) + ( Xd_0__inst_mult_0_37  ) + ( Xd_0__inst_mult_0_36  ))
// Xd_0__inst_mult_3_36  = CARRY(( (din_a[43] & din_b[36]) ) + ( Xd_0__inst_mult_0_37  ) + ( Xd_0__inst_mult_0_36  ))
// Xd_0__inst_mult_3_37  = SHARE(GND)

	.dataa(!din_a[43]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_36 ),
	.sharein(Xd_0__inst_mult_0_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_35_sumout ),
	.cout(Xd_0__inst_mult_3_36 ),
	.shareout(Xd_0__inst_mult_3_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_90 (
// Equation(s):
// Xd_0__inst_mult_9_272  = SUM(( (din_a[117] & din_b[112]) ) + ( Xd_0__inst_mult_9_386  ) + ( Xd_0__inst_mult_9_385  ))
// Xd_0__inst_mult_9_273  = CARRY(( (din_a[117] & din_b[112]) ) + ( Xd_0__inst_mult_9_386  ) + ( Xd_0__inst_mult_9_385  ))
// Xd_0__inst_mult_9_274  = SHARE(GND)

	.dataa(!din_a[117]),
	.datab(!din_b[112]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_385 ),
	.sharein(Xd_0__inst_mult_9_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_272 ),
	.cout(Xd_0__inst_mult_9_273 ),
	.shareout(Xd_0__inst_mult_9_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_91 (
// Equation(s):
// Xd_0__inst_mult_9_276  = SUM(( !Xd_0__inst_mult_9_388  $ (!Xd_0__inst_mult_9_384  $ (((din_b[110] & din_a[118])))) ) + ( Xd_0__inst_mult_9_342  ) + ( Xd_0__inst_mult_9_341  ))
// Xd_0__inst_mult_9_277  = CARRY(( !Xd_0__inst_mult_9_388  $ (!Xd_0__inst_mult_9_384  $ (((din_b[110] & din_a[118])))) ) + ( Xd_0__inst_mult_9_342  ) + ( Xd_0__inst_mult_9_341  ))
// Xd_0__inst_mult_9_278  = SHARE((!Xd_0__inst_mult_9_388  & (Xd_0__inst_mult_9_384  & (din_b[110] & din_a[118]))) # (Xd_0__inst_mult_9_388  & (((din_b[110] & din_a[118])) # (Xd_0__inst_mult_9_384 ))))

	.dataa(!Xd_0__inst_mult_9_388 ),
	.datab(!Xd_0__inst_mult_9_384 ),
	.datac(!din_b[110]),
	.datad(!din_a[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_341 ),
	.sharein(Xd_0__inst_mult_9_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_276 ),
	.cout(Xd_0__inst_mult_9_277 ),
	.shareout(Xd_0__inst_mult_9_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_43 (
// Equation(s):
// Xd_0__inst_mult_14_43_sumout  = SUM(( (din_a[178] & din_b[174]) ) + ( Xd_0__inst_mult_15_49  ) + ( Xd_0__inst_mult_15_48  ))
// Xd_0__inst_mult_14_44  = CARRY(( (din_a[178] & din_b[174]) ) + ( Xd_0__inst_mult_15_49  ) + ( Xd_0__inst_mult_15_48  ))
// Xd_0__inst_mult_14_45  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[174]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_48 ),
	.sharein(Xd_0__inst_mult_15_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_43_sumout ),
	.cout(Xd_0__inst_mult_14_44 ),
	.shareout(Xd_0__inst_mult_14_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_90 (
// Equation(s):
// Xd_0__inst_mult_6_272  = SUM(( (din_a[81] & din_b[76]) ) + ( Xd_0__inst_mult_6_386  ) + ( Xd_0__inst_mult_6_385  ))
// Xd_0__inst_mult_6_273  = CARRY(( (din_a[81] & din_b[76]) ) + ( Xd_0__inst_mult_6_386  ) + ( Xd_0__inst_mult_6_385  ))
// Xd_0__inst_mult_6_274  = SHARE(GND)

	.dataa(!din_a[81]),
	.datab(!din_b[76]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_385 ),
	.sharein(Xd_0__inst_mult_6_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_272 ),
	.cout(Xd_0__inst_mult_6_273 ),
	.shareout(Xd_0__inst_mult_6_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_91 (
// Equation(s):
// Xd_0__inst_mult_6_276  = SUM(( !Xd_0__inst_mult_6_388  $ (!Xd_0__inst_mult_6_384  $ (((din_b[74] & din_a[82])))) ) + ( Xd_0__inst_mult_6_342  ) + ( Xd_0__inst_mult_6_341  ))
// Xd_0__inst_mult_6_277  = CARRY(( !Xd_0__inst_mult_6_388  $ (!Xd_0__inst_mult_6_384  $ (((din_b[74] & din_a[82])))) ) + ( Xd_0__inst_mult_6_342  ) + ( Xd_0__inst_mult_6_341  ))
// Xd_0__inst_mult_6_278  = SHARE((!Xd_0__inst_mult_6_388  & (Xd_0__inst_mult_6_384  & (din_b[74] & din_a[82]))) # (Xd_0__inst_mult_6_388  & (((din_b[74] & din_a[82])) # (Xd_0__inst_mult_6_384 ))))

	.dataa(!Xd_0__inst_mult_6_388 ),
	.datab(!Xd_0__inst_mult_6_384 ),
	.datac(!din_b[74]),
	.datad(!din_a[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_341 ),
	.sharein(Xd_0__inst_mult_6_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_276 ),
	.cout(Xd_0__inst_mult_6_277 ),
	.shareout(Xd_0__inst_mult_6_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_99 (
// Equation(s):
// Xd_0__inst_mult_14_296  = SUM(( (!din_a[176] & (((din_a[175] & din_b[172])))) # (din_a[176] & (!din_b[171] $ (((!din_a[175]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_406  ) + ( Xd_0__inst_mult_14_405  ))
// Xd_0__inst_mult_14_297  = CARRY(( (!din_a[176] & (((din_a[175] & din_b[172])))) # (din_a[176] & (!din_b[171] $ (((!din_a[175]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_406  ) + ( Xd_0__inst_mult_14_405  ))
// Xd_0__inst_mult_14_298  = SHARE((din_a[176] & (din_b[171] & (din_a[175] & din_b[172]))))

	.dataa(!din_a[176]),
	.datab(!din_b[171]),
	.datac(!din_a[175]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_405 ),
	.sharein(Xd_0__inst_mult_14_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_296 ),
	.cout(Xd_0__inst_mult_14_297 ),
	.shareout(Xd_0__inst_mult_14_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_100 (
// Equation(s):
// Xd_0__inst_mult_14_300  = SUM(( (din_a[177] & din_b[170]) ) + ( Xd_0__inst_mult_14_410  ) + ( Xd_0__inst_mult_14_409  ))
// Xd_0__inst_mult_14_301  = CARRY(( (din_a[177] & din_b[170]) ) + ( Xd_0__inst_mult_14_410  ) + ( Xd_0__inst_mult_14_409  ))
// Xd_0__inst_mult_14_302  = SHARE(GND)

	.dataa(!din_a[177]),
	.datab(!din_b[170]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_409 ),
	.sharein(Xd_0__inst_mult_14_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_300 ),
	.cout(Xd_0__inst_mult_14_301 ),
	.shareout(Xd_0__inst_mult_14_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_101 (
// Equation(s):
// Xd_0__inst_mult_14_304  = SUM(( !Xd_0__inst_mult_14_408  $ (!Xd_0__inst_mult_14_404  $ (Xd_0__inst_mult_14_47_sumout )) ) + ( Xd_0__inst_mult_14_354  ) + ( Xd_0__inst_mult_14_353  ))
// Xd_0__inst_mult_14_305  = CARRY(( !Xd_0__inst_mult_14_408  $ (!Xd_0__inst_mult_14_404  $ (Xd_0__inst_mult_14_47_sumout )) ) + ( Xd_0__inst_mult_14_354  ) + ( Xd_0__inst_mult_14_353  ))
// Xd_0__inst_mult_14_306  = SHARE((!Xd_0__inst_mult_14_408  & (Xd_0__inst_mult_14_404  & Xd_0__inst_mult_14_47_sumout )) # (Xd_0__inst_mult_14_408  & ((Xd_0__inst_mult_14_47_sumout ) # (Xd_0__inst_mult_14_404 ))))

	.dataa(!Xd_0__inst_mult_14_408 ),
	.datab(!Xd_0__inst_mult_14_404 ),
	.datac(!Xd_0__inst_mult_14_47_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_353 ),
	.sharein(Xd_0__inst_mult_14_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_304 ),
	.cout(Xd_0__inst_mult_14_305 ),
	.shareout(Xd_0__inst_mult_14_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_94 (
// Equation(s):
// Xd_0__inst_mult_8_276  = SUM(( (din_a[105] & din_b[100]) ) + ( Xd_0__inst_mult_8_390  ) + ( Xd_0__inst_mult_8_389  ))
// Xd_0__inst_mult_8_277  = CARRY(( (din_a[105] & din_b[100]) ) + ( Xd_0__inst_mult_8_390  ) + ( Xd_0__inst_mult_8_389  ))
// Xd_0__inst_mult_8_278  = SHARE(GND)

	.dataa(!din_a[105]),
	.datab(!din_b[100]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_389 ),
	.sharein(Xd_0__inst_mult_8_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_276 ),
	.cout(Xd_0__inst_mult_8_277 ),
	.shareout(Xd_0__inst_mult_8_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_95 (
// Equation(s):
// Xd_0__inst_mult_8_280  = SUM(( !Xd_0__inst_mult_8_392  $ (!Xd_0__inst_mult_8_388  $ (((din_b[98] & din_a[106])))) ) + ( Xd_0__inst_mult_8_346  ) + ( Xd_0__inst_mult_8_345  ))
// Xd_0__inst_mult_8_281  = CARRY(( !Xd_0__inst_mult_8_392  $ (!Xd_0__inst_mult_8_388  $ (((din_b[98] & din_a[106])))) ) + ( Xd_0__inst_mult_8_346  ) + ( Xd_0__inst_mult_8_345  ))
// Xd_0__inst_mult_8_282  = SHARE((!Xd_0__inst_mult_8_392  & (Xd_0__inst_mult_8_388  & (din_b[98] & din_a[106]))) # (Xd_0__inst_mult_8_392  & (((din_b[98] & din_a[106])) # (Xd_0__inst_mult_8_388 ))))

	.dataa(!Xd_0__inst_mult_8_392 ),
	.datab(!Xd_0__inst_mult_8_388 ),
	.datac(!din_b[98]),
	.datad(!din_a[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_345 ),
	.sharein(Xd_0__inst_mult_8_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_280 ),
	.cout(Xd_0__inst_mult_8_281 ),
	.shareout(Xd_0__inst_mult_8_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_35 (
// Equation(s):
// Xd_0__inst_mult_9_35_sumout  = SUM(( (din_a[118] & din_b[115]) ) + ( Xd_0__inst_i29_23  ) + ( Xd_0__inst_i29_22  ))
// Xd_0__inst_mult_9_36  = CARRY(( (din_a[118] & din_b[115]) ) + ( Xd_0__inst_i29_23  ) + ( Xd_0__inst_i29_22  ))
// Xd_0__inst_mult_9_37  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[115]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_22 ),
	.sharein(Xd_0__inst_i29_23 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_35_sumout ),
	.cout(Xd_0__inst_mult_9_36 ),
	.shareout(Xd_0__inst_mult_9_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_94 (
// Equation(s):
// Xd_0__inst_mult_11_276  = SUM(( (din_a[141] & din_b[136]) ) + ( Xd_0__inst_mult_11_390  ) + ( Xd_0__inst_mult_11_389  ))
// Xd_0__inst_mult_11_277  = CARRY(( (din_a[141] & din_b[136]) ) + ( Xd_0__inst_mult_11_390  ) + ( Xd_0__inst_mult_11_389  ))
// Xd_0__inst_mult_11_278  = SHARE(GND)

	.dataa(!din_a[141]),
	.datab(!din_b[136]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_389 ),
	.sharein(Xd_0__inst_mult_11_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_276 ),
	.cout(Xd_0__inst_mult_11_277 ),
	.shareout(Xd_0__inst_mult_11_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_95 (
// Equation(s):
// Xd_0__inst_mult_11_280  = SUM(( !Xd_0__inst_mult_11_392  $ (!Xd_0__inst_mult_11_388  $ (((din_b[134] & din_a[142])))) ) + ( Xd_0__inst_mult_11_346  ) + ( Xd_0__inst_mult_11_345  ))
// Xd_0__inst_mult_11_281  = CARRY(( !Xd_0__inst_mult_11_392  $ (!Xd_0__inst_mult_11_388  $ (((din_b[134] & din_a[142])))) ) + ( Xd_0__inst_mult_11_346  ) + ( Xd_0__inst_mult_11_345  ))
// Xd_0__inst_mult_11_282  = SHARE((!Xd_0__inst_mult_11_392  & (Xd_0__inst_mult_11_388  & (din_b[134] & din_a[142]))) # (Xd_0__inst_mult_11_392  & (((din_b[134] & din_a[142])) # (Xd_0__inst_mult_11_388 ))))

	.dataa(!Xd_0__inst_mult_11_392 ),
	.datab(!Xd_0__inst_mult_11_388 ),
	.datac(!din_b[134]),
	.datad(!din_a[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_345 ),
	.sharein(Xd_0__inst_mult_11_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_280 ),
	.cout(Xd_0__inst_mult_11_281 ),
	.shareout(Xd_0__inst_mult_11_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_90 (
// Equation(s):
// Xd_0__inst_mult_10_272  = SUM(( (din_a[129] & din_b[124]) ) + ( Xd_0__inst_mult_10_386  ) + ( Xd_0__inst_mult_10_385  ))
// Xd_0__inst_mult_10_273  = CARRY(( (din_a[129] & din_b[124]) ) + ( Xd_0__inst_mult_10_386  ) + ( Xd_0__inst_mult_10_385  ))
// Xd_0__inst_mult_10_274  = SHARE(GND)

	.dataa(!din_a[129]),
	.datab(!din_b[124]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_385 ),
	.sharein(Xd_0__inst_mult_10_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_272 ),
	.cout(Xd_0__inst_mult_10_273 ),
	.shareout(Xd_0__inst_mult_10_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_91 (
// Equation(s):
// Xd_0__inst_mult_10_276  = SUM(( !Xd_0__inst_mult_10_388  $ (!Xd_0__inst_mult_10_384  $ (((din_b[122] & din_a[130])))) ) + ( Xd_0__inst_mult_10_342  ) + ( Xd_0__inst_mult_10_341  ))
// Xd_0__inst_mult_10_277  = CARRY(( !Xd_0__inst_mult_10_388  $ (!Xd_0__inst_mult_10_384  $ (((din_b[122] & din_a[130])))) ) + ( Xd_0__inst_mult_10_342  ) + ( Xd_0__inst_mult_10_341  ))
// Xd_0__inst_mult_10_278  = SHARE((!Xd_0__inst_mult_10_388  & (Xd_0__inst_mult_10_384  & (din_b[122] & din_a[130]))) # (Xd_0__inst_mult_10_388  & (((din_b[122] & din_a[130])) # (Xd_0__inst_mult_10_384 ))))

	.dataa(!Xd_0__inst_mult_10_388 ),
	.datab(!Xd_0__inst_mult_10_384 ),
	.datac(!din_b[122]),
	.datad(!din_a[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_341 ),
	.sharein(Xd_0__inst_mult_10_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_276 ),
	.cout(Xd_0__inst_mult_10_277 ),
	.shareout(Xd_0__inst_mult_10_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_99 (
// Equation(s):
// Xd_0__inst_mult_15_296  = SUM(( (din_a[185] & din_b[189]) ) + ( Xd_0__inst_mult_15_414  ) + ( Xd_0__inst_mult_15_413  ))
// Xd_0__inst_mult_15_297  = CARRY(( (din_a[185] & din_b[189]) ) + ( Xd_0__inst_mult_15_414  ) + ( Xd_0__inst_mult_15_413  ))
// Xd_0__inst_mult_15_298  = SHARE((din_a[185] & din_b[190]))

	.dataa(!din_a[185]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_413 ),
	.sharein(Xd_0__inst_mult_15_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_296 ),
	.cout(Xd_0__inst_mult_15_297 ),
	.shareout(Xd_0__inst_mult_15_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_94 (
// Equation(s):
// Xd_0__inst_mult_13_276  = SUM(( (din_a[165] & din_b[160]) ) + ( Xd_0__inst_mult_13_390  ) + ( Xd_0__inst_mult_13_389  ))
// Xd_0__inst_mult_13_277  = CARRY(( (din_a[165] & din_b[160]) ) + ( Xd_0__inst_mult_13_390  ) + ( Xd_0__inst_mult_13_389  ))
// Xd_0__inst_mult_13_278  = SHARE(GND)

	.dataa(!din_a[165]),
	.datab(!din_b[160]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_389 ),
	.sharein(Xd_0__inst_mult_13_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_276 ),
	.cout(Xd_0__inst_mult_13_277 ),
	.shareout(Xd_0__inst_mult_13_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_95 (
// Equation(s):
// Xd_0__inst_mult_13_280  = SUM(( !Xd_0__inst_mult_13_392  $ (!Xd_0__inst_mult_13_388  $ (((din_b[158] & din_a[166])))) ) + ( Xd_0__inst_mult_13_346  ) + ( Xd_0__inst_mult_13_345  ))
// Xd_0__inst_mult_13_281  = CARRY(( !Xd_0__inst_mult_13_392  $ (!Xd_0__inst_mult_13_388  $ (((din_b[158] & din_a[166])))) ) + ( Xd_0__inst_mult_13_346  ) + ( Xd_0__inst_mult_13_345  ))
// Xd_0__inst_mult_13_282  = SHARE((!Xd_0__inst_mult_13_392  & (Xd_0__inst_mult_13_388  & (din_b[158] & din_a[166]))) # (Xd_0__inst_mult_13_392  & (((din_b[158] & din_a[166])) # (Xd_0__inst_mult_13_388 ))))

	.dataa(!Xd_0__inst_mult_13_392 ),
	.datab(!Xd_0__inst_mult_13_388 ),
	.datac(!din_b[158]),
	.datad(!din_a[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_345 ),
	.sharein(Xd_0__inst_mult_13_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_280 ),
	.cout(Xd_0__inst_mult_13_281 ),
	.shareout(Xd_0__inst_mult_13_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_100 (
// Equation(s):
// Xd_0__inst_mult_15_300  = SUM(( (din_a[189] & din_b[184]) ) + ( Xd_0__inst_mult_15_418  ) + ( Xd_0__inst_mult_15_417  ))
// Xd_0__inst_mult_15_301  = CARRY(( (din_a[189] & din_b[184]) ) + ( Xd_0__inst_mult_15_418  ) + ( Xd_0__inst_mult_15_417  ))
// Xd_0__inst_mult_15_302  = SHARE(GND)

	.dataa(!din_a[189]),
	.datab(!din_b[184]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_417 ),
	.sharein(Xd_0__inst_mult_15_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_300 ),
	.cout(Xd_0__inst_mult_15_301 ),
	.shareout(Xd_0__inst_mult_15_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_101 (
// Equation(s):
// Xd_0__inst_mult_15_304  = SUM(( !Xd_0__inst_mult_15_420  $ (!Xd_0__inst_mult_15_416  $ (((din_b[182] & din_a[190])))) ) + ( Xd_0__inst_mult_15_370  ) + ( Xd_0__inst_mult_15_369  ))
// Xd_0__inst_mult_15_305  = CARRY(( !Xd_0__inst_mult_15_420  $ (!Xd_0__inst_mult_15_416  $ (((din_b[182] & din_a[190])))) ) + ( Xd_0__inst_mult_15_370  ) + ( Xd_0__inst_mult_15_369  ))
// Xd_0__inst_mult_15_306  = SHARE((!Xd_0__inst_mult_15_420  & (Xd_0__inst_mult_15_416  & (din_b[182] & din_a[190]))) # (Xd_0__inst_mult_15_420  & (((din_b[182] & din_a[190])) # (Xd_0__inst_mult_15_416 ))))

	.dataa(!Xd_0__inst_mult_15_420 ),
	.datab(!Xd_0__inst_mult_15_416 ),
	.datac(!din_b[182]),
	.datad(!din_a[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_369 ),
	.sharein(Xd_0__inst_mult_15_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_304 ),
	.cout(Xd_0__inst_mult_15_305 ),
	.shareout(Xd_0__inst_mult_15_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_95 (
// Equation(s):
// Xd_0__inst_mult_12_292  = SUM(( (din_a[153] & din_b[148]) ) + ( Xd_0__inst_mult_12_410  ) + ( Xd_0__inst_mult_12_409  ))
// Xd_0__inst_mult_12_293  = CARRY(( (din_a[153] & din_b[148]) ) + ( Xd_0__inst_mult_12_410  ) + ( Xd_0__inst_mult_12_409  ))
// Xd_0__inst_mult_12_294  = SHARE(GND)

	.dataa(!din_a[153]),
	.datab(!din_b[148]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_409 ),
	.sharein(Xd_0__inst_mult_12_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_292 ),
	.cout(Xd_0__inst_mult_12_293 ),
	.shareout(Xd_0__inst_mult_12_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_96 (
// Equation(s):
// Xd_0__inst_mult_12_296  = SUM(( !Xd_0__inst_mult_12_412  $ (!Xd_0__inst_mult_12_408  $ (((din_b[146] & din_a[154])))) ) + ( Xd_0__inst_mult_12_366  ) + ( Xd_0__inst_mult_12_365  ))
// Xd_0__inst_mult_12_297  = CARRY(( !Xd_0__inst_mult_12_412  $ (!Xd_0__inst_mult_12_408  $ (((din_b[146] & din_a[154])))) ) + ( Xd_0__inst_mult_12_366  ) + ( Xd_0__inst_mult_12_365  ))
// Xd_0__inst_mult_12_298  = SHARE((!Xd_0__inst_mult_12_412  & (Xd_0__inst_mult_12_408  & (din_b[146] & din_a[154]))) # (Xd_0__inst_mult_12_412  & (((din_b[146] & din_a[154])) # (Xd_0__inst_mult_12_408 ))))

	.dataa(!Xd_0__inst_mult_12_412 ),
	.datab(!Xd_0__inst_mult_12_408 ),
	.datac(!din_b[146]),
	.datad(!din_a[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_365 ),
	.sharein(Xd_0__inst_mult_12_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_296 ),
	.cout(Xd_0__inst_mult_12_297 ),
	.shareout(Xd_0__inst_mult_12_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_97 (
// Equation(s):
// Xd_0__inst_mult_12_300  = SUM(( (din_a[149] & din_b[153]) ) + ( Xd_0__inst_mult_12_418  ) + ( Xd_0__inst_mult_12_417  ))
// Xd_0__inst_mult_12_301  = CARRY(( (din_a[149] & din_b[153]) ) + ( Xd_0__inst_mult_12_418  ) + ( Xd_0__inst_mult_12_417  ))
// Xd_0__inst_mult_12_302  = SHARE((din_a[149] & din_b[154]))

	.dataa(!din_a[149]),
	.datab(!din_b[153]),
	.datac(!din_b[154]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_417 ),
	.sharein(Xd_0__inst_mult_12_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_300 ),
	.cout(Xd_0__inst_mult_12_301 ),
	.shareout(Xd_0__inst_mult_12_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_97 (
// Equation(s):
// Xd_0__inst_mult_4_288  = SUM(( (din_a[51] & din_b[57]) ) + ( Xd_0__inst_mult_4_414  ) + ( Xd_0__inst_mult_4_413  ))
// Xd_0__inst_mult_4_289  = CARRY(( (din_a[51] & din_b[57]) ) + ( Xd_0__inst_mult_4_414  ) + ( Xd_0__inst_mult_4_413  ))
// Xd_0__inst_mult_4_290  = SHARE((din_a[51] & din_b[58]))

	.dataa(!din_a[51]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_413 ),
	.sharein(Xd_0__inst_mult_4_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_288 ),
	.cout(Xd_0__inst_mult_4_289 ),
	.shareout(Xd_0__inst_mult_4_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_12_98 (
// Equation(s):
// Xd_0__inst_mult_12_305  = CARRY(( Xd_0__inst_mult_12_420  ) + ( Xd_0__inst_mult_12_426  ) + ( Xd_0__inst_mult_12_425  ))
// Xd_0__inst_mult_12_306  = SHARE((din_a[145] & din_b[146]))

	.dataa(!Xd_0__inst_mult_12_420 ),
	.datab(!din_a[145]),
	.datac(!din_b[146]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_425 ),
	.sharein(Xd_0__inst_mult_12_426 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_305 ),
	.shareout(Xd_0__inst_mult_12_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_13_96 (
// Equation(s):
// Xd_0__inst_mult_13_285  = CARRY(( Xd_0__inst_mult_13_396  ) + ( Xd_0__inst_mult_13_402  ) + ( Xd_0__inst_mult_13_401  ))
// Xd_0__inst_mult_13_286  = SHARE((din_a[157] & din_b[158]))

	.dataa(!Xd_0__inst_mult_13_396 ),
	.datab(!din_a[157]),
	.datac(!din_b[158]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_401 ),
	.sharein(Xd_0__inst_mult_13_402 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_285 ),
	.shareout(Xd_0__inst_mult_13_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_14_102 (
// Equation(s):
// Xd_0__inst_mult_14_309  = CARRY(( Xd_0__inst_mult_14_412  ) + ( Xd_0__inst_mult_14_418  ) + ( Xd_0__inst_mult_14_417  ))
// Xd_0__inst_mult_14_310  = SHARE((din_a[169] & din_b[170]))

	.dataa(!Xd_0__inst_mult_14_412 ),
	.datab(!din_a[169]),
	.datac(!din_b[170]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_417 ),
	.sharein(Xd_0__inst_mult_14_418 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_309 ),
	.shareout(Xd_0__inst_mult_14_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_15_102 (
// Equation(s):
// Xd_0__inst_mult_15_309  = CARRY(( Xd_0__inst_mult_15_424  ) + ( Xd_0__inst_mult_15_430  ) + ( Xd_0__inst_mult_15_429  ))
// Xd_0__inst_mult_15_310  = SHARE((din_a[181] & din_b[182]))

	.dataa(!Xd_0__inst_mult_15_424 ),
	.datab(!din_a[181]),
	.datac(!din_b[182]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_429 ),
	.sharein(Xd_0__inst_mult_15_430 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_309 ),
	.shareout(Xd_0__inst_mult_15_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_10_92 (
// Equation(s):
// Xd_0__inst_mult_10_281  = CARRY(( Xd_0__inst_mult_10_392  ) + ( Xd_0__inst_mult_10_398  ) + ( Xd_0__inst_mult_10_397  ))
// Xd_0__inst_mult_10_282  = SHARE((din_a[121] & din_b[122]))

	.dataa(!Xd_0__inst_mult_10_392 ),
	.datab(!din_a[121]),
	.datac(!din_b[122]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_397 ),
	.sharein(Xd_0__inst_mult_10_398 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_281 ),
	.shareout(Xd_0__inst_mult_10_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_11_96 (
// Equation(s):
// Xd_0__inst_mult_11_285  = CARRY(( Xd_0__inst_mult_11_396  ) + ( Xd_0__inst_mult_11_402  ) + ( Xd_0__inst_mult_11_401  ))
// Xd_0__inst_mult_11_286  = SHARE((din_a[133] & din_b[134]))

	.dataa(!Xd_0__inst_mult_11_396 ),
	.datab(!din_a[133]),
	.datac(!din_b[134]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_401 ),
	.sharein(Xd_0__inst_mult_11_402 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_285 ),
	.shareout(Xd_0__inst_mult_11_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_8_96 (
// Equation(s):
// Xd_0__inst_mult_8_285  = CARRY(( Xd_0__inst_mult_8_396  ) + ( Xd_0__inst_mult_8_402  ) + ( Xd_0__inst_mult_8_401  ))
// Xd_0__inst_mult_8_286  = SHARE((din_a[97] & din_b[98]))

	.dataa(!Xd_0__inst_mult_8_396 ),
	.datab(!din_a[97]),
	.datac(!din_b[98]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_401 ),
	.sharein(Xd_0__inst_mult_8_402 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_285 ),
	.shareout(Xd_0__inst_mult_8_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_9_92 (
// Equation(s):
// Xd_0__inst_mult_9_281  = CARRY(( Xd_0__inst_mult_9_392  ) + ( Xd_0__inst_mult_9_398  ) + ( Xd_0__inst_mult_9_397  ))
// Xd_0__inst_mult_9_282  = SHARE((din_a[109] & din_b[110]))

	.dataa(!Xd_0__inst_mult_9_392 ),
	.datab(!din_a[109]),
	.datac(!din_b[110]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_397 ),
	.sharein(Xd_0__inst_mult_9_398 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_281 ),
	.shareout(Xd_0__inst_mult_9_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_6_92 (
// Equation(s):
// Xd_0__inst_mult_6_281  = CARRY(( Xd_0__inst_mult_6_392  ) + ( Xd_0__inst_mult_6_398  ) + ( Xd_0__inst_mult_6_397  ))
// Xd_0__inst_mult_6_282  = SHARE((din_a[73] & din_b[74]))

	.dataa(!Xd_0__inst_mult_6_392 ),
	.datab(!din_a[73]),
	.datac(!din_b[74]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_397 ),
	.sharein(Xd_0__inst_mult_6_398 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_281 ),
	.shareout(Xd_0__inst_mult_6_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_7_86 (
// Equation(s):
// Xd_0__inst_mult_7_257  = CARRY(( Xd_0__inst_mult_7_376  ) + ( Xd_0__inst_mult_7_382  ) + ( Xd_0__inst_mult_7_381  ))
// Xd_0__inst_mult_7_258  = SHARE((din_a[85] & din_b[86]))

	.dataa(!Xd_0__inst_mult_7_376 ),
	.datab(!din_a[85]),
	.datac(!din_b[86]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_381 ),
	.sharein(Xd_0__inst_mult_7_382 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_257 ),
	.shareout(Xd_0__inst_mult_7_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_4_98 (
// Equation(s):
// Xd_0__inst_mult_4_293  = CARRY(( Xd_0__inst_mult_4_416  ) + ( Xd_0__inst_mult_4_422  ) + ( Xd_0__inst_mult_4_421  ))
// Xd_0__inst_mult_4_294  = SHARE((din_a[49] & din_b[50]))

	.dataa(!Xd_0__inst_mult_4_416 ),
	.datab(!din_a[49]),
	.datac(!din_b[50]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_421 ),
	.sharein(Xd_0__inst_mult_4_422 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_293 ),
	.shareout(Xd_0__inst_mult_4_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_5_86 (
// Equation(s):
// Xd_0__inst_mult_5_257  = CARRY(( Xd_0__inst_mult_5_376  ) + ( Xd_0__inst_mult_5_382  ) + ( Xd_0__inst_mult_5_381  ))
// Xd_0__inst_mult_5_258  = SHARE((din_a[61] & din_b[62]))

	.dataa(!Xd_0__inst_mult_5_376 ),
	.datab(!din_a[61]),
	.datac(!din_b[62]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_381 ),
	.sharein(Xd_0__inst_mult_5_382 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_257 ),
	.shareout(Xd_0__inst_mult_5_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_2_90 (
// Equation(s):
// Xd_0__inst_mult_2_261  = CARRY(( Xd_0__inst_mult_2_380  ) + ( Xd_0__inst_mult_2_386  ) + ( Xd_0__inst_mult_2_385  ))
// Xd_0__inst_mult_2_262  = SHARE((din_a[25] & din_b[26]))

	.dataa(!Xd_0__inst_mult_2_380 ),
	.datab(!din_a[25]),
	.datac(!din_b[26]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_385 ),
	.sharein(Xd_0__inst_mult_2_386 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_261 ),
	.shareout(Xd_0__inst_mult_2_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_3_86 (
// Equation(s):
// Xd_0__inst_mult_3_257  = CARRY(( Xd_0__inst_mult_3_376  ) + ( Xd_0__inst_mult_3_382  ) + ( Xd_0__inst_mult_3_381  ))
// Xd_0__inst_mult_3_258  = SHARE((din_a[37] & din_b[38]))

	.dataa(!Xd_0__inst_mult_3_376 ),
	.datab(!din_a[37]),
	.datac(!din_b[38]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_381 ),
	.sharein(Xd_0__inst_mult_3_382 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_257 ),
	.shareout(Xd_0__inst_mult_3_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_0_90 (
// Equation(s):
// Xd_0__inst_mult_0_261  = CARRY(( Xd_0__inst_mult_0_384  ) + ( Xd_0__inst_mult_0_362  ) + ( Xd_0__inst_mult_0_361  ))
// Xd_0__inst_mult_0_262  = SHARE((din_a[1] & din_b[2]))

	.dataa(!Xd_0__inst_mult_0_384 ),
	.datab(!din_a[1]),
	.datac(!din_b[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_361 ),
	.sharein(Xd_0__inst_mult_0_362 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_261 ),
	.shareout(Xd_0__inst_mult_0_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_1_90 (
// Equation(s):
// Xd_0__inst_mult_1_261  = CARRY(( Xd_0__inst_mult_1_384  ) + ( Xd_0__inst_mult_1_362  ) + ( Xd_0__inst_mult_1_361  ))
// Xd_0__inst_mult_1_262  = SHARE((din_a[13] & din_b[14]))

	.dataa(!Xd_0__inst_mult_1_384 ),
	.datab(!din_a[13]),
	.datac(!din_b[14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_361 ),
	.sharein(Xd_0__inst_mult_1_362 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_261 ),
	.shareout(Xd_0__inst_mult_1_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_99 (
// Equation(s):
// Xd_0__inst_mult_12_308  = SUM(( (din_a[148] & din_b[144]) ) + ( Xd_0__inst_mult_12_422  ) + ( Xd_0__inst_mult_12_421  ))
// Xd_0__inst_mult_12_309  = CARRY(( (din_a[148] & din_b[144]) ) + ( Xd_0__inst_mult_12_422  ) + ( Xd_0__inst_mult_12_421  ))
// Xd_0__inst_mult_12_310  = SHARE((din_a[148] & din_b[145]))

	.dataa(!din_a[148]),
	.datab(!din_b[144]),
	.datac(!din_b[145]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_421 ),
	.sharein(Xd_0__inst_mult_12_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_308 ),
	.cout(Xd_0__inst_mult_12_309 ),
	.shareout(Xd_0__inst_mult_12_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_100 (
// Equation(s):
// Xd_0__inst_mult_12_312  = SUM(( (din_a[145] & din_b[147]) ) + ( Xd_0__inst_mult_12_430  ) + ( Xd_0__inst_mult_12_429  ))
// Xd_0__inst_mult_12_313  = CARRY(( (din_a[145] & din_b[147]) ) + ( Xd_0__inst_mult_12_430  ) + ( Xd_0__inst_mult_12_429  ))
// Xd_0__inst_mult_12_314  = SHARE((din_b[147] & din_a[146]))

	.dataa(!din_a[145]),
	.datab(!din_b[147]),
	.datac(!din_a[146]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_429 ),
	.sharein(Xd_0__inst_mult_12_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_312 ),
	.cout(Xd_0__inst_mult_12_313 ),
	.shareout(Xd_0__inst_mult_12_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_97 (
// Equation(s):
// Xd_0__inst_mult_13_288  = SUM(( (din_a[160] & din_b[156]) ) + ( Xd_0__inst_mult_13_398  ) + ( Xd_0__inst_mult_13_397  ))
// Xd_0__inst_mult_13_289  = CARRY(( (din_a[160] & din_b[156]) ) + ( Xd_0__inst_mult_13_398  ) + ( Xd_0__inst_mult_13_397  ))
// Xd_0__inst_mult_13_290  = SHARE((din_a[160] & din_b[157]))

	.dataa(!din_a[160]),
	.datab(!din_b[156]),
	.datac(!din_b[157]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_397 ),
	.sharein(Xd_0__inst_mult_13_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_288 ),
	.cout(Xd_0__inst_mult_13_289 ),
	.shareout(Xd_0__inst_mult_13_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_98 (
// Equation(s):
// Xd_0__inst_mult_13_292  = SUM(( (din_a[157] & din_b[159]) ) + ( Xd_0__inst_mult_13_406  ) + ( Xd_0__inst_mult_13_405  ))
// Xd_0__inst_mult_13_293  = CARRY(( (din_a[157] & din_b[159]) ) + ( Xd_0__inst_mult_13_406  ) + ( Xd_0__inst_mult_13_405  ))
// Xd_0__inst_mult_13_294  = SHARE((din_b[159] & din_a[158]))

	.dataa(!din_a[157]),
	.datab(!din_b[159]),
	.datac(!din_a[158]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_405 ),
	.sharein(Xd_0__inst_mult_13_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_292 ),
	.cout(Xd_0__inst_mult_13_293 ),
	.shareout(Xd_0__inst_mult_13_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_103 (
// Equation(s):
// Xd_0__inst_mult_14_312  = SUM(( (din_a[172] & din_b[168]) ) + ( Xd_0__inst_mult_14_414  ) + ( Xd_0__inst_mult_14_413  ))
// Xd_0__inst_mult_14_313  = CARRY(( (din_a[172] & din_b[168]) ) + ( Xd_0__inst_mult_14_414  ) + ( Xd_0__inst_mult_14_413  ))
// Xd_0__inst_mult_14_314  = SHARE((din_a[172] & din_b[169]))

	.dataa(!din_a[172]),
	.datab(!din_b[168]),
	.datac(!din_b[169]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_413 ),
	.sharein(Xd_0__inst_mult_14_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_312 ),
	.cout(Xd_0__inst_mult_14_313 ),
	.shareout(Xd_0__inst_mult_14_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_104 (
// Equation(s):
// Xd_0__inst_mult_14_316  = SUM(( (din_a[169] & din_b[171]) ) + ( Xd_0__inst_mult_14_422  ) + ( Xd_0__inst_mult_14_421  ))
// Xd_0__inst_mult_14_317  = CARRY(( (din_a[169] & din_b[171]) ) + ( Xd_0__inst_mult_14_422  ) + ( Xd_0__inst_mult_14_421  ))
// Xd_0__inst_mult_14_318  = SHARE((din_b[171] & din_a[170]))

	.dataa(!din_a[169]),
	.datab(!din_b[171]),
	.datac(!din_a[170]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_421 ),
	.sharein(Xd_0__inst_mult_14_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_316 ),
	.cout(Xd_0__inst_mult_14_317 ),
	.shareout(Xd_0__inst_mult_14_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_103 (
// Equation(s):
// Xd_0__inst_mult_15_312  = SUM(( (din_a[184] & din_b[180]) ) + ( Xd_0__inst_mult_15_426  ) + ( Xd_0__inst_mult_15_425  ))
// Xd_0__inst_mult_15_313  = CARRY(( (din_a[184] & din_b[180]) ) + ( Xd_0__inst_mult_15_426  ) + ( Xd_0__inst_mult_15_425  ))
// Xd_0__inst_mult_15_314  = SHARE((din_a[184] & din_b[181]))

	.dataa(!din_a[184]),
	.datab(!din_b[180]),
	.datac(!din_b[181]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_425 ),
	.sharein(Xd_0__inst_mult_15_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_312 ),
	.cout(Xd_0__inst_mult_15_313 ),
	.shareout(Xd_0__inst_mult_15_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_104 (
// Equation(s):
// Xd_0__inst_mult_15_316  = SUM(( (din_a[181] & din_b[183]) ) + ( Xd_0__inst_mult_15_434  ) + ( Xd_0__inst_mult_15_433  ))
// Xd_0__inst_mult_15_317  = CARRY(( (din_a[181] & din_b[183]) ) + ( Xd_0__inst_mult_15_434  ) + ( Xd_0__inst_mult_15_433  ))
// Xd_0__inst_mult_15_318  = SHARE((din_b[183] & din_a[182]))

	.dataa(!din_a[181]),
	.datab(!din_b[183]),
	.datac(!din_a[182]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_433 ),
	.sharein(Xd_0__inst_mult_15_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_316 ),
	.cout(Xd_0__inst_mult_15_317 ),
	.shareout(Xd_0__inst_mult_15_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_93 (
// Equation(s):
// Xd_0__inst_mult_10_284  = SUM(( (din_a[124] & din_b[120]) ) + ( Xd_0__inst_mult_10_394  ) + ( Xd_0__inst_mult_10_393  ))
// Xd_0__inst_mult_10_285  = CARRY(( (din_a[124] & din_b[120]) ) + ( Xd_0__inst_mult_10_394  ) + ( Xd_0__inst_mult_10_393  ))
// Xd_0__inst_mult_10_286  = SHARE((din_a[124] & din_b[121]))

	.dataa(!din_a[124]),
	.datab(!din_b[120]),
	.datac(!din_b[121]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_393 ),
	.sharein(Xd_0__inst_mult_10_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_284 ),
	.cout(Xd_0__inst_mult_10_285 ),
	.shareout(Xd_0__inst_mult_10_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_94 (
// Equation(s):
// Xd_0__inst_mult_10_288  = SUM(( (din_a[121] & din_b[123]) ) + ( Xd_0__inst_mult_10_402  ) + ( Xd_0__inst_mult_10_401  ))
// Xd_0__inst_mult_10_289  = CARRY(( (din_a[121] & din_b[123]) ) + ( Xd_0__inst_mult_10_402  ) + ( Xd_0__inst_mult_10_401  ))
// Xd_0__inst_mult_10_290  = SHARE((din_b[123] & din_a[122]))

	.dataa(!din_a[121]),
	.datab(!din_b[123]),
	.datac(!din_a[122]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_401 ),
	.sharein(Xd_0__inst_mult_10_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_288 ),
	.cout(Xd_0__inst_mult_10_289 ),
	.shareout(Xd_0__inst_mult_10_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_97 (
// Equation(s):
// Xd_0__inst_mult_11_288  = SUM(( (din_a[136] & din_b[132]) ) + ( Xd_0__inst_mult_11_398  ) + ( Xd_0__inst_mult_11_397  ))
// Xd_0__inst_mult_11_289  = CARRY(( (din_a[136] & din_b[132]) ) + ( Xd_0__inst_mult_11_398  ) + ( Xd_0__inst_mult_11_397  ))
// Xd_0__inst_mult_11_290  = SHARE((din_a[136] & din_b[133]))

	.dataa(!din_a[136]),
	.datab(!din_b[132]),
	.datac(!din_b[133]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_397 ),
	.sharein(Xd_0__inst_mult_11_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_288 ),
	.cout(Xd_0__inst_mult_11_289 ),
	.shareout(Xd_0__inst_mult_11_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_98 (
// Equation(s):
// Xd_0__inst_mult_11_292  = SUM(( (din_a[133] & din_b[135]) ) + ( Xd_0__inst_mult_11_406  ) + ( Xd_0__inst_mult_11_405  ))
// Xd_0__inst_mult_11_293  = CARRY(( (din_a[133] & din_b[135]) ) + ( Xd_0__inst_mult_11_406  ) + ( Xd_0__inst_mult_11_405  ))
// Xd_0__inst_mult_11_294  = SHARE((din_b[135] & din_a[134]))

	.dataa(!din_a[133]),
	.datab(!din_b[135]),
	.datac(!din_a[134]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_405 ),
	.sharein(Xd_0__inst_mult_11_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_292 ),
	.cout(Xd_0__inst_mult_11_293 ),
	.shareout(Xd_0__inst_mult_11_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_97 (
// Equation(s):
// Xd_0__inst_mult_8_288  = SUM(( (din_a[100] & din_b[96]) ) + ( Xd_0__inst_mult_8_398  ) + ( Xd_0__inst_mult_8_397  ))
// Xd_0__inst_mult_8_289  = CARRY(( (din_a[100] & din_b[96]) ) + ( Xd_0__inst_mult_8_398  ) + ( Xd_0__inst_mult_8_397  ))
// Xd_0__inst_mult_8_290  = SHARE((din_a[100] & din_b[97]))

	.dataa(!din_a[100]),
	.datab(!din_b[96]),
	.datac(!din_b[97]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_397 ),
	.sharein(Xd_0__inst_mult_8_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_288 ),
	.cout(Xd_0__inst_mult_8_289 ),
	.shareout(Xd_0__inst_mult_8_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_98 (
// Equation(s):
// Xd_0__inst_mult_8_292  = SUM(( (din_a[97] & din_b[99]) ) + ( Xd_0__inst_mult_8_406  ) + ( Xd_0__inst_mult_8_405  ))
// Xd_0__inst_mult_8_293  = CARRY(( (din_a[97] & din_b[99]) ) + ( Xd_0__inst_mult_8_406  ) + ( Xd_0__inst_mult_8_405  ))
// Xd_0__inst_mult_8_294  = SHARE((din_b[99] & din_a[98]))

	.dataa(!din_a[97]),
	.datab(!din_b[99]),
	.datac(!din_a[98]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_405 ),
	.sharein(Xd_0__inst_mult_8_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_292 ),
	.cout(Xd_0__inst_mult_8_293 ),
	.shareout(Xd_0__inst_mult_8_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_93 (
// Equation(s):
// Xd_0__inst_mult_9_284  = SUM(( (din_a[112] & din_b[108]) ) + ( Xd_0__inst_mult_9_394  ) + ( Xd_0__inst_mult_9_393  ))
// Xd_0__inst_mult_9_285  = CARRY(( (din_a[112] & din_b[108]) ) + ( Xd_0__inst_mult_9_394  ) + ( Xd_0__inst_mult_9_393  ))
// Xd_0__inst_mult_9_286  = SHARE((din_a[112] & din_b[109]))

	.dataa(!din_a[112]),
	.datab(!din_b[108]),
	.datac(!din_b[109]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_393 ),
	.sharein(Xd_0__inst_mult_9_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_284 ),
	.cout(Xd_0__inst_mult_9_285 ),
	.shareout(Xd_0__inst_mult_9_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_94 (
// Equation(s):
// Xd_0__inst_mult_9_288  = SUM(( (din_a[109] & din_b[111]) ) + ( Xd_0__inst_mult_9_402  ) + ( Xd_0__inst_mult_9_401  ))
// Xd_0__inst_mult_9_289  = CARRY(( (din_a[109] & din_b[111]) ) + ( Xd_0__inst_mult_9_402  ) + ( Xd_0__inst_mult_9_401  ))
// Xd_0__inst_mult_9_290  = SHARE((din_b[111] & din_a[110]))

	.dataa(!din_a[109]),
	.datab(!din_b[111]),
	.datac(!din_a[110]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_401 ),
	.sharein(Xd_0__inst_mult_9_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_288 ),
	.cout(Xd_0__inst_mult_9_289 ),
	.shareout(Xd_0__inst_mult_9_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_93 (
// Equation(s):
// Xd_0__inst_mult_6_284  = SUM(( (din_a[76] & din_b[72]) ) + ( Xd_0__inst_mult_6_394  ) + ( Xd_0__inst_mult_6_393  ))
// Xd_0__inst_mult_6_285  = CARRY(( (din_a[76] & din_b[72]) ) + ( Xd_0__inst_mult_6_394  ) + ( Xd_0__inst_mult_6_393  ))
// Xd_0__inst_mult_6_286  = SHARE((din_a[76] & din_b[73]))

	.dataa(!din_a[76]),
	.datab(!din_b[72]),
	.datac(!din_b[73]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_393 ),
	.sharein(Xd_0__inst_mult_6_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_284 ),
	.cout(Xd_0__inst_mult_6_285 ),
	.shareout(Xd_0__inst_mult_6_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_94 (
// Equation(s):
// Xd_0__inst_mult_6_288  = SUM(( (din_a[73] & din_b[75]) ) + ( Xd_0__inst_mult_6_402  ) + ( Xd_0__inst_mult_6_401  ))
// Xd_0__inst_mult_6_289  = CARRY(( (din_a[73] & din_b[75]) ) + ( Xd_0__inst_mult_6_402  ) + ( Xd_0__inst_mult_6_401  ))
// Xd_0__inst_mult_6_290  = SHARE((din_b[75] & din_a[74]))

	.dataa(!din_a[73]),
	.datab(!din_b[75]),
	.datac(!din_a[74]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_401 ),
	.sharein(Xd_0__inst_mult_6_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_288 ),
	.cout(Xd_0__inst_mult_6_289 ),
	.shareout(Xd_0__inst_mult_6_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_87 (
// Equation(s):
// Xd_0__inst_mult_7_260  = SUM(( (din_a[88] & din_b[84]) ) + ( Xd_0__inst_mult_7_378  ) + ( Xd_0__inst_mult_7_377  ))
// Xd_0__inst_mult_7_261  = CARRY(( (din_a[88] & din_b[84]) ) + ( Xd_0__inst_mult_7_378  ) + ( Xd_0__inst_mult_7_377  ))
// Xd_0__inst_mult_7_262  = SHARE((din_a[88] & din_b[85]))

	.dataa(!din_a[88]),
	.datab(!din_b[84]),
	.datac(!din_b[85]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_377 ),
	.sharein(Xd_0__inst_mult_7_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_260 ),
	.cout(Xd_0__inst_mult_7_261 ),
	.shareout(Xd_0__inst_mult_7_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_88 (
// Equation(s):
// Xd_0__inst_mult_7_264  = SUM(( (din_a[85] & din_b[87]) ) + ( Xd_0__inst_mult_7_386  ) + ( Xd_0__inst_mult_7_385  ))
// Xd_0__inst_mult_7_265  = CARRY(( (din_a[85] & din_b[87]) ) + ( Xd_0__inst_mult_7_386  ) + ( Xd_0__inst_mult_7_385  ))
// Xd_0__inst_mult_7_266  = SHARE((din_b[87] & din_a[86]))

	.dataa(!din_a[85]),
	.datab(!din_b[87]),
	.datac(!din_a[86]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_385 ),
	.sharein(Xd_0__inst_mult_7_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_264 ),
	.cout(Xd_0__inst_mult_7_265 ),
	.shareout(Xd_0__inst_mult_7_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_99 (
// Equation(s):
// Xd_0__inst_mult_4_296  = SUM(( (din_a[52] & din_b[48]) ) + ( Xd_0__inst_mult_4_418  ) + ( Xd_0__inst_mult_4_417  ))
// Xd_0__inst_mult_4_297  = CARRY(( (din_a[52] & din_b[48]) ) + ( Xd_0__inst_mult_4_418  ) + ( Xd_0__inst_mult_4_417  ))
// Xd_0__inst_mult_4_298  = SHARE((din_a[52] & din_b[49]))

	.dataa(!din_a[52]),
	.datab(!din_b[48]),
	.datac(!din_b[49]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_417 ),
	.sharein(Xd_0__inst_mult_4_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_296 ),
	.cout(Xd_0__inst_mult_4_297 ),
	.shareout(Xd_0__inst_mult_4_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_100 (
// Equation(s):
// Xd_0__inst_mult_4_300  = SUM(( (din_a[49] & din_b[51]) ) + ( Xd_0__inst_mult_4_426  ) + ( Xd_0__inst_mult_4_425  ))
// Xd_0__inst_mult_4_301  = CARRY(( (din_a[49] & din_b[51]) ) + ( Xd_0__inst_mult_4_426  ) + ( Xd_0__inst_mult_4_425  ))
// Xd_0__inst_mult_4_302  = SHARE((din_b[51] & din_a[50]))

	.dataa(!din_a[49]),
	.datab(!din_b[51]),
	.datac(!din_a[50]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_425 ),
	.sharein(Xd_0__inst_mult_4_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_300 ),
	.cout(Xd_0__inst_mult_4_301 ),
	.shareout(Xd_0__inst_mult_4_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_87 (
// Equation(s):
// Xd_0__inst_mult_5_260  = SUM(( (din_a[64] & din_b[60]) ) + ( Xd_0__inst_mult_5_378  ) + ( Xd_0__inst_mult_5_377  ))
// Xd_0__inst_mult_5_261  = CARRY(( (din_a[64] & din_b[60]) ) + ( Xd_0__inst_mult_5_378  ) + ( Xd_0__inst_mult_5_377  ))
// Xd_0__inst_mult_5_262  = SHARE((din_a[64] & din_b[61]))

	.dataa(!din_a[64]),
	.datab(!din_b[60]),
	.datac(!din_b[61]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_377 ),
	.sharein(Xd_0__inst_mult_5_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_260 ),
	.cout(Xd_0__inst_mult_5_261 ),
	.shareout(Xd_0__inst_mult_5_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_88 (
// Equation(s):
// Xd_0__inst_mult_5_264  = SUM(( (din_a[61] & din_b[63]) ) + ( Xd_0__inst_mult_5_386  ) + ( Xd_0__inst_mult_5_385  ))
// Xd_0__inst_mult_5_265  = CARRY(( (din_a[61] & din_b[63]) ) + ( Xd_0__inst_mult_5_386  ) + ( Xd_0__inst_mult_5_385  ))
// Xd_0__inst_mult_5_266  = SHARE((din_b[63] & din_a[62]))

	.dataa(!din_a[61]),
	.datab(!din_b[63]),
	.datac(!din_a[62]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_385 ),
	.sharein(Xd_0__inst_mult_5_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_264 ),
	.cout(Xd_0__inst_mult_5_265 ),
	.shareout(Xd_0__inst_mult_5_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_91 (
// Equation(s):
// Xd_0__inst_mult_2_264  = SUM(( (din_a[28] & din_b[24]) ) + ( Xd_0__inst_mult_2_382  ) + ( Xd_0__inst_mult_2_381  ))
// Xd_0__inst_mult_2_265  = CARRY(( (din_a[28] & din_b[24]) ) + ( Xd_0__inst_mult_2_382  ) + ( Xd_0__inst_mult_2_381  ))
// Xd_0__inst_mult_2_266  = SHARE((din_a[28] & din_b[25]))

	.dataa(!din_a[28]),
	.datab(!din_b[24]),
	.datac(!din_b[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_381 ),
	.sharein(Xd_0__inst_mult_2_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_264 ),
	.cout(Xd_0__inst_mult_2_265 ),
	.shareout(Xd_0__inst_mult_2_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_92 (
// Equation(s):
// Xd_0__inst_mult_2_268  = SUM(( (din_a[25] & din_b[27]) ) + ( Xd_0__inst_mult_2_390  ) + ( Xd_0__inst_mult_2_389  ))
// Xd_0__inst_mult_2_269  = CARRY(( (din_a[25] & din_b[27]) ) + ( Xd_0__inst_mult_2_390  ) + ( Xd_0__inst_mult_2_389  ))
// Xd_0__inst_mult_2_270  = SHARE((din_b[27] & din_a[26]))

	.dataa(!din_a[25]),
	.datab(!din_b[27]),
	.datac(!din_a[26]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_389 ),
	.sharein(Xd_0__inst_mult_2_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_268 ),
	.cout(Xd_0__inst_mult_2_269 ),
	.shareout(Xd_0__inst_mult_2_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_87 (
// Equation(s):
// Xd_0__inst_mult_3_260  = SUM(( (din_a[40] & din_b[36]) ) + ( Xd_0__inst_mult_3_378  ) + ( Xd_0__inst_mult_3_377  ))
// Xd_0__inst_mult_3_261  = CARRY(( (din_a[40] & din_b[36]) ) + ( Xd_0__inst_mult_3_378  ) + ( Xd_0__inst_mult_3_377  ))
// Xd_0__inst_mult_3_262  = SHARE((din_a[40] & din_b[37]))

	.dataa(!din_a[40]),
	.datab(!din_b[36]),
	.datac(!din_b[37]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_377 ),
	.sharein(Xd_0__inst_mult_3_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_260 ),
	.cout(Xd_0__inst_mult_3_261 ),
	.shareout(Xd_0__inst_mult_3_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_88 (
// Equation(s):
// Xd_0__inst_mult_3_264  = SUM(( (din_a[37] & din_b[39]) ) + ( Xd_0__inst_mult_3_386  ) + ( Xd_0__inst_mult_3_385  ))
// Xd_0__inst_mult_3_265  = CARRY(( (din_a[37] & din_b[39]) ) + ( Xd_0__inst_mult_3_386  ) + ( Xd_0__inst_mult_3_385  ))
// Xd_0__inst_mult_3_266  = SHARE((din_b[39] & din_a[38]))

	.dataa(!din_a[37]),
	.datab(!din_b[39]),
	.datac(!din_a[38]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_385 ),
	.sharein(Xd_0__inst_mult_3_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_264 ),
	.cout(Xd_0__inst_mult_3_265 ),
	.shareout(Xd_0__inst_mult_3_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_91 (
// Equation(s):
// Xd_0__inst_mult_0_264  = SUM(( (din_a[4] & din_b[0]) ) + ( Xd_0__inst_mult_0_386  ) + ( Xd_0__inst_mult_0_385  ))
// Xd_0__inst_mult_0_265  = CARRY(( (din_a[4] & din_b[0]) ) + ( Xd_0__inst_mult_0_386  ) + ( Xd_0__inst_mult_0_385  ))
// Xd_0__inst_mult_0_266  = SHARE((din_a[4] & din_b[1]))

	.dataa(!din_a[4]),
	.datab(!din_b[0]),
	.datac(!din_b[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_385 ),
	.sharein(Xd_0__inst_mult_0_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_264 ),
	.cout(Xd_0__inst_mult_0_265 ),
	.shareout(Xd_0__inst_mult_0_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_92 (
// Equation(s):
// Xd_0__inst_mult_0_268  = SUM(( (din_a[1] & din_b[3]) ) + ( Xd_0__inst_mult_0_390  ) + ( Xd_0__inst_mult_0_389  ))
// Xd_0__inst_mult_0_269  = CARRY(( (din_a[1] & din_b[3]) ) + ( Xd_0__inst_mult_0_390  ) + ( Xd_0__inst_mult_0_389  ))
// Xd_0__inst_mult_0_270  = SHARE((din_b[3] & din_a[2]))

	.dataa(!din_a[1]),
	.datab(!din_b[3]),
	.datac(!din_a[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_389 ),
	.sharein(Xd_0__inst_mult_0_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_268 ),
	.cout(Xd_0__inst_mult_0_269 ),
	.shareout(Xd_0__inst_mult_0_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_91 (
// Equation(s):
// Xd_0__inst_mult_1_264  = SUM(( (din_a[16] & din_b[12]) ) + ( Xd_0__inst_mult_1_386  ) + ( Xd_0__inst_mult_1_385  ))
// Xd_0__inst_mult_1_265  = CARRY(( (din_a[16] & din_b[12]) ) + ( Xd_0__inst_mult_1_386  ) + ( Xd_0__inst_mult_1_385  ))
// Xd_0__inst_mult_1_266  = SHARE((din_a[16] & din_b[13]))

	.dataa(!din_a[16]),
	.datab(!din_b[12]),
	.datac(!din_b[13]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_385 ),
	.sharein(Xd_0__inst_mult_1_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_264 ),
	.cout(Xd_0__inst_mult_1_265 ),
	.shareout(Xd_0__inst_mult_1_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_92 (
// Equation(s):
// Xd_0__inst_mult_1_268  = SUM(( (din_a[13] & din_b[15]) ) + ( Xd_0__inst_mult_1_390  ) + ( Xd_0__inst_mult_1_389  ))
// Xd_0__inst_mult_1_269  = CARRY(( (din_a[13] & din_b[15]) ) + ( Xd_0__inst_mult_1_390  ) + ( Xd_0__inst_mult_1_389  ))
// Xd_0__inst_mult_1_270  = SHARE((din_b[15] & din_a[14]))

	.dataa(!din_a[13]),
	.datab(!din_b[15]),
	.datac(!din_a[14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_389 ),
	.sharein(Xd_0__inst_mult_1_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_268 ),
	.cout(Xd_0__inst_mult_1_269 ),
	.shareout(Xd_0__inst_mult_1_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_101 (
// Equation(s):
// Xd_0__inst_mult_12_316  = SUM(( !Xd_0__inst_mult_12_432  $ (!Xd_0__inst_mult_12_436  $ (((din_b[148] & din_a[145])))) ) + ( Xd_0__inst_mult_12_290  ) + ( Xd_0__inst_mult_12_289  ))
// Xd_0__inst_mult_12_317  = CARRY(( !Xd_0__inst_mult_12_432  $ (!Xd_0__inst_mult_12_436  $ (((din_b[148] & din_a[145])))) ) + ( Xd_0__inst_mult_12_290  ) + ( Xd_0__inst_mult_12_289  ))
// Xd_0__inst_mult_12_318  = SHARE((!Xd_0__inst_mult_12_432  & (Xd_0__inst_mult_12_436  & (din_b[148] & din_a[145]))) # (Xd_0__inst_mult_12_432  & (((din_b[148] & din_a[145])) # (Xd_0__inst_mult_12_436 ))))

	.dataa(!Xd_0__inst_mult_12_432 ),
	.datab(!Xd_0__inst_mult_12_436 ),
	.datac(!din_b[148]),
	.datad(!din_a[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_289 ),
	.sharein(Xd_0__inst_mult_12_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_316 ),
	.cout(Xd_0__inst_mult_12_317 ),
	.shareout(Xd_0__inst_mult_12_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_102 (
// Equation(s):
// Xd_0__inst_mult_12_320  = SUM(( (din_a[144] & din_b[149]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_321  = CARRY(( (din_a[144] & din_b[149]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_322  = SHARE((din_a[144] & din_b[150]))

	.dataa(!din_a[144]),
	.datab(!din_b[149]),
	.datac(!din_b[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_12_320 ),
	.cout(Xd_0__inst_mult_12_321 ),
	.shareout(Xd_0__inst_mult_12_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_39 (
// Equation(s):
// Xd_0__inst_mult_13_39_sumout  = SUM(( (din_a[166] & din_b[156]) ) + ( Xd_0__inst_mult_10_61  ) + ( Xd_0__inst_mult_10_60  ))
// Xd_0__inst_mult_13_40  = CARRY(( (din_a[166] & din_b[156]) ) + ( Xd_0__inst_mult_10_61  ) + ( Xd_0__inst_mult_10_60  ))
// Xd_0__inst_mult_13_41  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_60 ),
	.sharein(Xd_0__inst_mult_10_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_39_sumout ),
	.cout(Xd_0__inst_mult_13_40 ),
	.shareout(Xd_0__inst_mult_13_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_99 (
// Equation(s):
// Xd_0__inst_mult_13_296  = SUM(( !Xd_0__inst_mult_13_408  $ (!Xd_0__inst_mult_13_412  $ (((din_b[160] & din_a[157])))) ) + ( Xd_0__inst_mult_13_274  ) + ( Xd_0__inst_mult_13_273  ))
// Xd_0__inst_mult_13_297  = CARRY(( !Xd_0__inst_mult_13_408  $ (!Xd_0__inst_mult_13_412  $ (((din_b[160] & din_a[157])))) ) + ( Xd_0__inst_mult_13_274  ) + ( Xd_0__inst_mult_13_273  ))
// Xd_0__inst_mult_13_298  = SHARE((!Xd_0__inst_mult_13_408  & (Xd_0__inst_mult_13_412  & (din_b[160] & din_a[157]))) # (Xd_0__inst_mult_13_408  & (((din_b[160] & din_a[157])) # (Xd_0__inst_mult_13_412 ))))

	.dataa(!Xd_0__inst_mult_13_408 ),
	.datab(!Xd_0__inst_mult_13_412 ),
	.datac(!din_b[160]),
	.datad(!din_a[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_273 ),
	.sharein(Xd_0__inst_mult_13_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_296 ),
	.cout(Xd_0__inst_mult_13_297 ),
	.shareout(Xd_0__inst_mult_13_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_100 (
// Equation(s):
// Xd_0__inst_mult_13_300  = SUM(( (din_a[156] & din_b[161]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_301  = CARRY(( (din_a[156] & din_b[161]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_302  = SHARE((din_a[156] & din_b[162]))

	.dataa(!din_a[156]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_13_300 ),
	.cout(Xd_0__inst_mult_13_301 ),
	.shareout(Xd_0__inst_mult_13_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_47 (
// Equation(s):
// Xd_0__inst_mult_14_47_sumout  = SUM(( (din_a[178] & din_b[168]) ) + ( Xd_0__inst_mult_15_65  ) + ( Xd_0__inst_mult_15_64  ))
// Xd_0__inst_mult_14_48  = CARRY(( (din_a[178] & din_b[168]) ) + ( Xd_0__inst_mult_15_65  ) + ( Xd_0__inst_mult_15_64  ))
// Xd_0__inst_mult_14_49  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[168]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_64 ),
	.sharein(Xd_0__inst_mult_15_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_47_sumout ),
	.cout(Xd_0__inst_mult_14_48 ),
	.shareout(Xd_0__inst_mult_14_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_105 (
// Equation(s):
// Xd_0__inst_mult_14_320  = SUM(( !Xd_0__inst_mult_14_424  $ (!Xd_0__inst_mult_14_428  $ (((din_b[172] & din_a[169])))) ) + ( Xd_0__inst_mult_14_294  ) + ( Xd_0__inst_mult_14_293  ))
// Xd_0__inst_mult_14_321  = CARRY(( !Xd_0__inst_mult_14_424  $ (!Xd_0__inst_mult_14_428  $ (((din_b[172] & din_a[169])))) ) + ( Xd_0__inst_mult_14_294  ) + ( Xd_0__inst_mult_14_293  ))
// Xd_0__inst_mult_14_322  = SHARE((!Xd_0__inst_mult_14_424  & (Xd_0__inst_mult_14_428  & (din_b[172] & din_a[169]))) # (Xd_0__inst_mult_14_424  & (((din_b[172] & din_a[169])) # (Xd_0__inst_mult_14_428 ))))

	.dataa(!Xd_0__inst_mult_14_424 ),
	.datab(!Xd_0__inst_mult_14_428 ),
	.datac(!din_b[172]),
	.datad(!din_a[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_293 ),
	.sharein(Xd_0__inst_mult_14_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_320 ),
	.cout(Xd_0__inst_mult_14_321 ),
	.shareout(Xd_0__inst_mult_14_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_106 (
// Equation(s):
// Xd_0__inst_mult_14_324  = SUM(( (din_a[168] & din_b[173]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_325  = CARRY(( (din_a[168] & din_b[173]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_326  = SHARE((din_a[168] & din_b[174]))

	.dataa(!din_a[168]),
	.datab(!din_b[173]),
	.datac(!din_b[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_14_324 ),
	.cout(Xd_0__inst_mult_14_325 ),
	.shareout(Xd_0__inst_mult_14_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_35 (
// Equation(s):
// Xd_0__inst_mult_7_35_sumout  = SUM(( (din_a[94] & din_b[84]) ) + ( Xd_0__inst_mult_4_57  ) + ( Xd_0__inst_mult_4_56  ))
// Xd_0__inst_mult_7_36  = CARRY(( (din_a[94] & din_b[84]) ) + ( Xd_0__inst_mult_4_57  ) + ( Xd_0__inst_mult_4_56  ))
// Xd_0__inst_mult_7_37  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_56 ),
	.sharein(Xd_0__inst_mult_4_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_35_sumout ),
	.cout(Xd_0__inst_mult_7_36 ),
	.shareout(Xd_0__inst_mult_7_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_105 (
// Equation(s):
// Xd_0__inst_mult_15_320  = SUM(( !Xd_0__inst_mult_15_436  $ (!Xd_0__inst_mult_15_440  $ (((din_b[184] & din_a[181])))) ) + ( Xd_0__inst_mult_15_294  ) + ( Xd_0__inst_mult_15_293  ))
// Xd_0__inst_mult_15_321  = CARRY(( !Xd_0__inst_mult_15_436  $ (!Xd_0__inst_mult_15_440  $ (((din_b[184] & din_a[181])))) ) + ( Xd_0__inst_mult_15_294  ) + ( Xd_0__inst_mult_15_293  ))
// Xd_0__inst_mult_15_322  = SHARE((!Xd_0__inst_mult_15_436  & (Xd_0__inst_mult_15_440  & (din_b[184] & din_a[181]))) # (Xd_0__inst_mult_15_436  & (((din_b[184] & din_a[181])) # (Xd_0__inst_mult_15_440 ))))

	.dataa(!Xd_0__inst_mult_15_436 ),
	.datab(!Xd_0__inst_mult_15_440 ),
	.datac(!din_b[184]),
	.datad(!din_a[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_293 ),
	.sharein(Xd_0__inst_mult_15_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_320 ),
	.cout(Xd_0__inst_mult_15_321 ),
	.shareout(Xd_0__inst_mult_15_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_106 (
// Equation(s):
// Xd_0__inst_mult_15_324  = SUM(( (din_a[180] & din_b[185]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_325  = CARRY(( (din_a[180] & din_b[185]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_326  = SHARE((din_a[180] & din_b[186]))

	.dataa(!din_a[180]),
	.datab(!din_b[185]),
	.datac(!din_b[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_15_324 ),
	.cout(Xd_0__inst_mult_15_325 ),
	.shareout(Xd_0__inst_mult_15_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_35 (
// Equation(s):
// Xd_0__inst_mult_8_35_sumout  = SUM(( (din_a[106] & din_b[96]) ) + ( Xd_0__inst_mult_9_57  ) + ( Xd_0__inst_mult_9_56  ))
// Xd_0__inst_mult_8_36  = CARRY(( (din_a[106] & din_b[96]) ) + ( Xd_0__inst_mult_9_57  ) + ( Xd_0__inst_mult_9_56  ))
// Xd_0__inst_mult_8_37  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[96]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_56 ),
	.sharein(Xd_0__inst_mult_9_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_35_sumout ),
	.cout(Xd_0__inst_mult_8_36 ),
	.shareout(Xd_0__inst_mult_8_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_95 (
// Equation(s):
// Xd_0__inst_mult_10_292  = SUM(( !Xd_0__inst_mult_10_404  $ (!Xd_0__inst_mult_10_408  $ (((din_b[124] & din_a[121])))) ) + ( Xd_0__inst_mult_10_270  ) + ( Xd_0__inst_mult_10_269  ))
// Xd_0__inst_mult_10_293  = CARRY(( !Xd_0__inst_mult_10_404  $ (!Xd_0__inst_mult_10_408  $ (((din_b[124] & din_a[121])))) ) + ( Xd_0__inst_mult_10_270  ) + ( Xd_0__inst_mult_10_269  ))
// Xd_0__inst_mult_10_294  = SHARE((!Xd_0__inst_mult_10_404  & (Xd_0__inst_mult_10_408  & (din_b[124] & din_a[121]))) # (Xd_0__inst_mult_10_404  & (((din_b[124] & din_a[121])) # (Xd_0__inst_mult_10_408 ))))

	.dataa(!Xd_0__inst_mult_10_404 ),
	.datab(!Xd_0__inst_mult_10_408 ),
	.datac(!din_b[124]),
	.datad(!din_a[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_269 ),
	.sharein(Xd_0__inst_mult_10_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_292 ),
	.cout(Xd_0__inst_mult_10_293 ),
	.shareout(Xd_0__inst_mult_10_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_96 (
// Equation(s):
// Xd_0__inst_mult_10_296  = SUM(( (din_a[120] & din_b[125]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_297  = CARRY(( (din_a[120] & din_b[125]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_298  = SHARE((din_a[120] & din_b[126]))

	.dataa(!din_a[120]),
	.datab(!din_b[125]),
	.datac(!din_b[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_10_296 ),
	.cout(Xd_0__inst_mult_10_297 ),
	.shareout(Xd_0__inst_mult_10_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_39 (
// Equation(s):
// Xd_0__inst_mult_3_39_sumout  = SUM(( (din_a[45] & din_b[36]) ) + ( Xd_0__inst_mult_0_61  ) + ( Xd_0__inst_mult_0_60  ))
// Xd_0__inst_mult_3_40  = CARRY(( (din_a[45] & din_b[36]) ) + ( Xd_0__inst_mult_0_61  ) + ( Xd_0__inst_mult_0_60  ))
// Xd_0__inst_mult_3_41  = SHARE(GND)

	.dataa(!din_a[45]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_60 ),
	.sharein(Xd_0__inst_mult_0_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_39_sumout ),
	.cout(Xd_0__inst_mult_3_40 ),
	.shareout(Xd_0__inst_mult_3_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_99 (
// Equation(s):
// Xd_0__inst_mult_11_296  = SUM(( !Xd_0__inst_mult_11_408  $ (!Xd_0__inst_mult_11_412  $ (((din_b[136] & din_a[133])))) ) + ( Xd_0__inst_mult_11_274  ) + ( Xd_0__inst_mult_11_273  ))
// Xd_0__inst_mult_11_297  = CARRY(( !Xd_0__inst_mult_11_408  $ (!Xd_0__inst_mult_11_412  $ (((din_b[136] & din_a[133])))) ) + ( Xd_0__inst_mult_11_274  ) + ( Xd_0__inst_mult_11_273  ))
// Xd_0__inst_mult_11_298  = SHARE((!Xd_0__inst_mult_11_408  & (Xd_0__inst_mult_11_412  & (din_b[136] & din_a[133]))) # (Xd_0__inst_mult_11_408  & (((din_b[136] & din_a[133])) # (Xd_0__inst_mult_11_412 ))))

	.dataa(!Xd_0__inst_mult_11_408 ),
	.datab(!Xd_0__inst_mult_11_412 ),
	.datac(!din_b[136]),
	.datad(!din_a[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_273 ),
	.sharein(Xd_0__inst_mult_11_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_296 ),
	.cout(Xd_0__inst_mult_11_297 ),
	.shareout(Xd_0__inst_mult_11_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_100 (
// Equation(s):
// Xd_0__inst_mult_11_300  = SUM(( (din_a[132] & din_b[137]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_301  = CARRY(( (din_a[132] & din_b[137]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_302  = SHARE((din_a[132] & din_b[138]))

	.dataa(!din_a[132]),
	.datab(!din_b[137]),
	.datac(!din_b[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_300 ),
	.cout(Xd_0__inst_mult_11_301 ),
	.shareout(Xd_0__inst_mult_11_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_39 (
// Equation(s):
// Xd_0__inst_mult_15_39_sumout  = SUM(( (din_a[187] & din_b[180]) ) + ( Xd_0__inst_mult_11_57  ) + ( Xd_0__inst_mult_11_56  ))
// Xd_0__inst_mult_15_40  = CARRY(( (din_a[187] & din_b[180]) ) + ( Xd_0__inst_mult_11_57  ) + ( Xd_0__inst_mult_11_56  ))
// Xd_0__inst_mult_15_41  = SHARE(GND)

	.dataa(!din_a[187]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_56 ),
	.sharein(Xd_0__inst_mult_11_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_39_sumout ),
	.cout(Xd_0__inst_mult_15_40 ),
	.shareout(Xd_0__inst_mult_15_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_99 (
// Equation(s):
// Xd_0__inst_mult_8_296  = SUM(( !Xd_0__inst_mult_8_408  $ (!Xd_0__inst_mult_8_412  $ (((din_b[100] & din_a[97])))) ) + ( Xd_0__inst_mult_8_274  ) + ( Xd_0__inst_mult_8_273  ))
// Xd_0__inst_mult_8_297  = CARRY(( !Xd_0__inst_mult_8_408  $ (!Xd_0__inst_mult_8_412  $ (((din_b[100] & din_a[97])))) ) + ( Xd_0__inst_mult_8_274  ) + ( Xd_0__inst_mult_8_273  ))
// Xd_0__inst_mult_8_298  = SHARE((!Xd_0__inst_mult_8_408  & (Xd_0__inst_mult_8_412  & (din_b[100] & din_a[97]))) # (Xd_0__inst_mult_8_408  & (((din_b[100] & din_a[97])) # (Xd_0__inst_mult_8_412 ))))

	.dataa(!Xd_0__inst_mult_8_408 ),
	.datab(!Xd_0__inst_mult_8_412 ),
	.datac(!din_b[100]),
	.datad(!din_a[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_273 ),
	.sharein(Xd_0__inst_mult_8_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_296 ),
	.cout(Xd_0__inst_mult_8_297 ),
	.shareout(Xd_0__inst_mult_8_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_100 (
// Equation(s):
// Xd_0__inst_mult_8_300  = SUM(( (din_a[96] & din_b[101]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_301  = CARRY(( (din_a[96] & din_b[101]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_302  = SHARE((din_a[96] & din_b[102]))

	.dataa(!din_a[96]),
	.datab(!din_b[101]),
	.datac(!din_b[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_8_300 ),
	.cout(Xd_0__inst_mult_8_301 ),
	.shareout(Xd_0__inst_mult_8_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_43 (
// Equation(s):
// Xd_0__inst_mult_3_43_sumout  = SUM(( (din_a[46] & din_b[46]) ) + ( Xd_0__inst_mult_0_57  ) + ( Xd_0__inst_mult_0_56  ))
// Xd_0__inst_mult_3_44  = CARRY(( (din_a[46] & din_b[46]) ) + ( Xd_0__inst_mult_0_57  ) + ( Xd_0__inst_mult_0_56  ))
// Xd_0__inst_mult_3_45  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_56 ),
	.sharein(Xd_0__inst_mult_0_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_43_sumout ),
	.cout(Xd_0__inst_mult_3_44 ),
	.shareout(Xd_0__inst_mult_3_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_95 (
// Equation(s):
// Xd_0__inst_mult_9_292  = SUM(( !Xd_0__inst_mult_9_404  $ (!Xd_0__inst_mult_9_408  $ (((din_b[112] & din_a[109])))) ) + ( Xd_0__inst_mult_9_270  ) + ( Xd_0__inst_mult_9_269  ))
// Xd_0__inst_mult_9_293  = CARRY(( !Xd_0__inst_mult_9_404  $ (!Xd_0__inst_mult_9_408  $ (((din_b[112] & din_a[109])))) ) + ( Xd_0__inst_mult_9_270  ) + ( Xd_0__inst_mult_9_269  ))
// Xd_0__inst_mult_9_294  = SHARE((!Xd_0__inst_mult_9_404  & (Xd_0__inst_mult_9_408  & (din_b[112] & din_a[109]))) # (Xd_0__inst_mult_9_404  & (((din_b[112] & din_a[109])) # (Xd_0__inst_mult_9_408 ))))

	.dataa(!Xd_0__inst_mult_9_404 ),
	.datab(!Xd_0__inst_mult_9_408 ),
	.datac(!din_b[112]),
	.datad(!din_a[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_269 ),
	.sharein(Xd_0__inst_mult_9_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_292 ),
	.cout(Xd_0__inst_mult_9_293 ),
	.shareout(Xd_0__inst_mult_9_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_96 (
// Equation(s):
// Xd_0__inst_mult_9_296  = SUM(( (din_a[108] & din_b[113]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_297  = CARRY(( (din_a[108] & din_b[113]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_298  = SHARE((din_a[108] & din_b[114]))

	.dataa(!din_a[108]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_296 ),
	.cout(Xd_0__inst_mult_9_297 ),
	.shareout(Xd_0__inst_mult_9_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_39 (
// Equation(s):
// Xd_0__inst_mult_1_39_sumout  = SUM(( (din_a[22] & din_b[12]) ) + ( Xd_0__inst_mult_1_61  ) + ( Xd_0__inst_mult_1_60  ))
// Xd_0__inst_mult_1_40  = CARRY(( (din_a[22] & din_b[12]) ) + ( Xd_0__inst_mult_1_61  ) + ( Xd_0__inst_mult_1_60  ))
// Xd_0__inst_mult_1_41  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_60 ),
	.sharein(Xd_0__inst_mult_1_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_39_sumout ),
	.cout(Xd_0__inst_mult_1_40 ),
	.shareout(Xd_0__inst_mult_1_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_95 (
// Equation(s):
// Xd_0__inst_mult_6_292  = SUM(( !Xd_0__inst_mult_6_404  $ (!Xd_0__inst_mult_6_408  $ (((din_b[76] & din_a[73])))) ) + ( Xd_0__inst_mult_6_270  ) + ( Xd_0__inst_mult_6_269  ))
// Xd_0__inst_mult_6_293  = CARRY(( !Xd_0__inst_mult_6_404  $ (!Xd_0__inst_mult_6_408  $ (((din_b[76] & din_a[73])))) ) + ( Xd_0__inst_mult_6_270  ) + ( Xd_0__inst_mult_6_269  ))
// Xd_0__inst_mult_6_294  = SHARE((!Xd_0__inst_mult_6_404  & (Xd_0__inst_mult_6_408  & (din_b[76] & din_a[73]))) # (Xd_0__inst_mult_6_404  & (((din_b[76] & din_a[73])) # (Xd_0__inst_mult_6_408 ))))

	.dataa(!Xd_0__inst_mult_6_404 ),
	.datab(!Xd_0__inst_mult_6_408 ),
	.datac(!din_b[76]),
	.datad(!din_a[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_269 ),
	.sharein(Xd_0__inst_mult_6_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_292 ),
	.cout(Xd_0__inst_mult_6_293 ),
	.shareout(Xd_0__inst_mult_6_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_96 (
// Equation(s):
// Xd_0__inst_mult_6_296  = SUM(( (din_a[72] & din_b[77]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_297  = CARRY(( (din_a[72] & din_b[77]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_298  = SHARE((din_a[72] & din_b[78]))

	.dataa(!din_a[72]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_296 ),
	.cout(Xd_0__inst_mult_6_297 ),
	.shareout(Xd_0__inst_mult_6_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_43 (
// Equation(s):
// Xd_0__inst_mult_12_43_sumout  = SUM(( (din_a[151] & din_b[144]) ) + ( Xd_0__inst_mult_13_61  ) + ( Xd_0__inst_mult_13_60  ))
// Xd_0__inst_mult_12_44  = CARRY(( (din_a[151] & din_b[144]) ) + ( Xd_0__inst_mult_13_61  ) + ( Xd_0__inst_mult_13_60  ))
// Xd_0__inst_mult_12_45  = SHARE(GND)

	.dataa(!din_a[151]),
	.datab(!din_b[144]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_60 ),
	.sharein(Xd_0__inst_mult_13_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_43_sumout ),
	.cout(Xd_0__inst_mult_12_44 ),
	.shareout(Xd_0__inst_mult_12_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_89 (
// Equation(s):
// Xd_0__inst_mult_7_268  = SUM(( !Xd_0__inst_mult_7_388  $ (!Xd_0__inst_mult_7_392  $ (((din_b[88] & din_a[85])))) ) + ( Xd_0__inst_mult_7_254  ) + ( Xd_0__inst_mult_7_253  ))
// Xd_0__inst_mult_7_269  = CARRY(( !Xd_0__inst_mult_7_388  $ (!Xd_0__inst_mult_7_392  $ (((din_b[88] & din_a[85])))) ) + ( Xd_0__inst_mult_7_254  ) + ( Xd_0__inst_mult_7_253  ))
// Xd_0__inst_mult_7_270  = SHARE((!Xd_0__inst_mult_7_388  & (Xd_0__inst_mult_7_392  & (din_b[88] & din_a[85]))) # (Xd_0__inst_mult_7_388  & (((din_b[88] & din_a[85])) # (Xd_0__inst_mult_7_392 ))))

	.dataa(!Xd_0__inst_mult_7_388 ),
	.datab(!Xd_0__inst_mult_7_392 ),
	.datac(!din_b[88]),
	.datad(!din_a[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_253 ),
	.sharein(Xd_0__inst_mult_7_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_268 ),
	.cout(Xd_0__inst_mult_7_269 ),
	.shareout(Xd_0__inst_mult_7_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_90 (
// Equation(s):
// Xd_0__inst_mult_7_272  = SUM(( (din_a[84] & din_b[89]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_273  = CARRY(( (din_a[84] & din_b[89]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_274  = SHARE((din_a[84] & din_b[90]))

	.dataa(!din_a[84]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_272 ),
	.cout(Xd_0__inst_mult_7_273 ),
	.shareout(Xd_0__inst_mult_7_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_35 (
// Equation(s):
// Xd_0__inst_mult_11_35_sumout  = SUM(( (din_a[142] & din_b[142]) ) + ( Xd_0__inst_mult_10_57  ) + ( Xd_0__inst_mult_10_56  ))
// Xd_0__inst_mult_11_36  = CARRY(( (din_a[142] & din_b[142]) ) + ( Xd_0__inst_mult_10_57  ) + ( Xd_0__inst_mult_10_56  ))
// Xd_0__inst_mult_11_37  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_56 ),
	.sharein(Xd_0__inst_mult_10_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_35_sumout ),
	.cout(Xd_0__inst_mult_11_36 ),
	.shareout(Xd_0__inst_mult_11_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_101 (
// Equation(s):
// Xd_0__inst_mult_4_304  = SUM(( !Xd_0__inst_mult_4_428  $ (!Xd_0__inst_mult_4_432  $ (((din_b[52] & din_a[49])))) ) + ( Xd_0__inst_mult_4_286  ) + ( Xd_0__inst_mult_4_285  ))
// Xd_0__inst_mult_4_305  = CARRY(( !Xd_0__inst_mult_4_428  $ (!Xd_0__inst_mult_4_432  $ (((din_b[52] & din_a[49])))) ) + ( Xd_0__inst_mult_4_286  ) + ( Xd_0__inst_mult_4_285  ))
// Xd_0__inst_mult_4_306  = SHARE((!Xd_0__inst_mult_4_428  & (Xd_0__inst_mult_4_432  & (din_b[52] & din_a[49]))) # (Xd_0__inst_mult_4_428  & (((din_b[52] & din_a[49])) # (Xd_0__inst_mult_4_432 ))))

	.dataa(!Xd_0__inst_mult_4_428 ),
	.datab(!Xd_0__inst_mult_4_432 ),
	.datac(!din_b[52]),
	.datad(!din_a[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_285 ),
	.sharein(Xd_0__inst_mult_4_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_304 ),
	.cout(Xd_0__inst_mult_4_305 ),
	.shareout(Xd_0__inst_mult_4_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_102 (
// Equation(s):
// Xd_0__inst_mult_4_308  = SUM(( (din_a[48] & din_b[53]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_309  = CARRY(( (din_a[48] & din_b[53]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_310  = SHARE((din_a[48] & din_b[54]))

	.dataa(!din_a[48]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_308 ),
	.cout(Xd_0__inst_mult_4_309 ),
	.shareout(Xd_0__inst_mult_4_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_39 (
// Equation(s):
// Xd_0__inst_mult_8_39_sumout  = SUM(( (din_a[104] & din_b[96]) ) + ( Xd_0__inst_mult_2_61  ) + ( Xd_0__inst_mult_2_60  ))
// Xd_0__inst_mult_8_40  = CARRY(( (din_a[104] & din_b[96]) ) + ( Xd_0__inst_mult_2_61  ) + ( Xd_0__inst_mult_2_60  ))
// Xd_0__inst_mult_8_41  = SHARE(GND)

	.dataa(!din_a[104]),
	.datab(!din_b[96]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_60 ),
	.sharein(Xd_0__inst_mult_2_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_39_sumout ),
	.cout(Xd_0__inst_mult_8_40 ),
	.shareout(Xd_0__inst_mult_8_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_89 (
// Equation(s):
// Xd_0__inst_mult_5_268  = SUM(( !Xd_0__inst_mult_5_388  $ (!Xd_0__inst_mult_5_392  $ (((din_b[64] & din_a[61])))) ) + ( Xd_0__inst_mult_5_254  ) + ( Xd_0__inst_mult_5_253  ))
// Xd_0__inst_mult_5_269  = CARRY(( !Xd_0__inst_mult_5_388  $ (!Xd_0__inst_mult_5_392  $ (((din_b[64] & din_a[61])))) ) + ( Xd_0__inst_mult_5_254  ) + ( Xd_0__inst_mult_5_253  ))
// Xd_0__inst_mult_5_270  = SHARE((!Xd_0__inst_mult_5_388  & (Xd_0__inst_mult_5_392  & (din_b[64] & din_a[61]))) # (Xd_0__inst_mult_5_388  & (((din_b[64] & din_a[61])) # (Xd_0__inst_mult_5_392 ))))

	.dataa(!Xd_0__inst_mult_5_388 ),
	.datab(!Xd_0__inst_mult_5_392 ),
	.datac(!din_b[64]),
	.datad(!din_a[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_253 ),
	.sharein(Xd_0__inst_mult_5_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_268 ),
	.cout(Xd_0__inst_mult_5_269 ),
	.shareout(Xd_0__inst_mult_5_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_90 (
// Equation(s):
// Xd_0__inst_mult_5_272  = SUM(( (din_a[60] & din_b[65]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_273  = CARRY(( (din_a[60] & din_b[65]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_274  = SHARE((din_a[60] & din_b[66]))

	.dataa(!din_a[60]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_272 ),
	.cout(Xd_0__inst_mult_5_273 ),
	.shareout(Xd_0__inst_mult_5_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_43 (
// Equation(s):
// Xd_0__inst_mult_8_43_sumout  = SUM(( (din_a[106] & din_b[106]) ) + ( Xd_0__inst_mult_7_53  ) + ( Xd_0__inst_mult_7_52  ))
// Xd_0__inst_mult_8_44  = CARRY(( (din_a[106] & din_b[106]) ) + ( Xd_0__inst_mult_7_53  ) + ( Xd_0__inst_mult_7_52  ))
// Xd_0__inst_mult_8_45  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[106]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_52 ),
	.sharein(Xd_0__inst_mult_7_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_43_sumout ),
	.cout(Xd_0__inst_mult_8_44 ),
	.shareout(Xd_0__inst_mult_8_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_93 (
// Equation(s):
// Xd_0__inst_mult_2_272  = SUM(( !Xd_0__inst_mult_2_392  $ (!Xd_0__inst_mult_2_396  $ (((din_b[28] & din_a[25])))) ) + ( Xd_0__inst_mult_2_258  ) + ( Xd_0__inst_mult_2_257  ))
// Xd_0__inst_mult_2_273  = CARRY(( !Xd_0__inst_mult_2_392  $ (!Xd_0__inst_mult_2_396  $ (((din_b[28] & din_a[25])))) ) + ( Xd_0__inst_mult_2_258  ) + ( Xd_0__inst_mult_2_257  ))
// Xd_0__inst_mult_2_274  = SHARE((!Xd_0__inst_mult_2_392  & (Xd_0__inst_mult_2_396  & (din_b[28] & din_a[25]))) # (Xd_0__inst_mult_2_392  & (((din_b[28] & din_a[25])) # (Xd_0__inst_mult_2_396 ))))

	.dataa(!Xd_0__inst_mult_2_392 ),
	.datab(!Xd_0__inst_mult_2_396 ),
	.datac(!din_b[28]),
	.datad(!din_a[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_257 ),
	.sharein(Xd_0__inst_mult_2_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_272 ),
	.cout(Xd_0__inst_mult_2_273 ),
	.shareout(Xd_0__inst_mult_2_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_94 (
// Equation(s):
// Xd_0__inst_mult_2_276  = SUM(( (din_a[24] & din_b[29]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_277  = CARRY(( (din_a[24] & din_b[29]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_278  = SHARE((din_a[24] & din_b[30]))

	.dataa(!din_a[24]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_276 ),
	.cout(Xd_0__inst_mult_2_277 ),
	.shareout(Xd_0__inst_mult_2_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_51 (
// Equation(s):
// Xd_0__inst_mult_14_51_sumout  = SUM(( (din_a[178] & din_b[178]) ) + ( Xd_0__inst_mult_9_53  ) + ( Xd_0__inst_mult_9_52  ))
// Xd_0__inst_mult_14_52  = CARRY(( (din_a[178] & din_b[178]) ) + ( Xd_0__inst_mult_9_53  ) + ( Xd_0__inst_mult_9_52  ))
// Xd_0__inst_mult_14_53  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[178]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_52 ),
	.sharein(Xd_0__inst_mult_9_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_51_sumout ),
	.cout(Xd_0__inst_mult_14_52 ),
	.shareout(Xd_0__inst_mult_14_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_89 (
// Equation(s):
// Xd_0__inst_mult_3_268  = SUM(( !Xd_0__inst_mult_3_388  $ (!Xd_0__inst_mult_3_392  $ (((din_b[40] & din_a[37])))) ) + ( Xd_0__inst_mult_3_254  ) + ( Xd_0__inst_mult_3_253  ))
// Xd_0__inst_mult_3_269  = CARRY(( !Xd_0__inst_mult_3_388  $ (!Xd_0__inst_mult_3_392  $ (((din_b[40] & din_a[37])))) ) + ( Xd_0__inst_mult_3_254  ) + ( Xd_0__inst_mult_3_253  ))
// Xd_0__inst_mult_3_270  = SHARE((!Xd_0__inst_mult_3_388  & (Xd_0__inst_mult_3_392  & (din_b[40] & din_a[37]))) # (Xd_0__inst_mult_3_388  & (((din_b[40] & din_a[37])) # (Xd_0__inst_mult_3_392 ))))

	.dataa(!Xd_0__inst_mult_3_388 ),
	.datab(!Xd_0__inst_mult_3_392 ),
	.datac(!din_b[40]),
	.datad(!din_a[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_253 ),
	.sharein(Xd_0__inst_mult_3_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_268 ),
	.cout(Xd_0__inst_mult_3_269 ),
	.shareout(Xd_0__inst_mult_3_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_90 (
// Equation(s):
// Xd_0__inst_mult_3_272  = SUM(( (din_a[36] & din_b[41]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_273  = CARRY(( (din_a[36] & din_b[41]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_274  = SHARE((din_a[36] & din_b[42]))

	.dataa(!din_a[36]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_272 ),
	.cout(Xd_0__inst_mult_3_273 ),
	.shareout(Xd_0__inst_mult_3_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_39 (
// Equation(s):
// Xd_0__inst_mult_10_39_sumout  = SUM(( (din_a[128] & din_b[120]) ) + ( Xd_0__inst_mult_11_61  ) + ( Xd_0__inst_mult_11_60  ))
// Xd_0__inst_mult_10_40  = CARRY(( (din_a[128] & din_b[120]) ) + ( Xd_0__inst_mult_11_61  ) + ( Xd_0__inst_mult_11_60  ))
// Xd_0__inst_mult_10_41  = SHARE(GND)

	.dataa(!din_a[128]),
	.datab(!din_b[120]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_60 ),
	.sharein(Xd_0__inst_mult_11_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_39_sumout ),
	.cout(Xd_0__inst_mult_10_40 ),
	.shareout(Xd_0__inst_mult_10_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_93 (
// Equation(s):
// Xd_0__inst_mult_0_272  = SUM(( !Xd_0__inst_mult_0_392  $ (!Xd_0__inst_mult_0_396  $ (((din_b[4] & din_a[1])))) ) + ( Xd_0__inst_mult_0_258  ) + ( Xd_0__inst_mult_0_257  ))
// Xd_0__inst_mult_0_273  = CARRY(( !Xd_0__inst_mult_0_392  $ (!Xd_0__inst_mult_0_396  $ (((din_b[4] & din_a[1])))) ) + ( Xd_0__inst_mult_0_258  ) + ( Xd_0__inst_mult_0_257  ))
// Xd_0__inst_mult_0_274  = SHARE((!Xd_0__inst_mult_0_392  & (Xd_0__inst_mult_0_396  & (din_b[4] & din_a[1]))) # (Xd_0__inst_mult_0_392  & (((din_b[4] & din_a[1])) # (Xd_0__inst_mult_0_396 ))))

	.dataa(!Xd_0__inst_mult_0_392 ),
	.datab(!Xd_0__inst_mult_0_396 ),
	.datac(!din_b[4]),
	.datad(!din_a[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_257 ),
	.sharein(Xd_0__inst_mult_0_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_272 ),
	.cout(Xd_0__inst_mult_0_273 ),
	.shareout(Xd_0__inst_mult_0_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_94 (
// Equation(s):
// Xd_0__inst_mult_0_276  = SUM(( (din_a[0] & din_b[5]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_277  = CARRY(( (din_a[0] & din_b[5]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_278  = SHARE((din_a[0] & din_b[6]))

	.dataa(!din_a[0]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_276 ),
	.cout(Xd_0__inst_mult_0_277 ),
	.shareout(Xd_0__inst_mult_0_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_43 (
// Equation(s):
// Xd_0__inst_mult_15_43_sumout  = SUM(( (din_a[188] & din_b[180]) ) + ( Xd_0__inst_mult_12_65  ) + ( Xd_0__inst_mult_12_64  ))
// Xd_0__inst_mult_15_44  = CARRY(( (din_a[188] & din_b[180]) ) + ( Xd_0__inst_mult_12_65  ) + ( Xd_0__inst_mult_12_64  ))
// Xd_0__inst_mult_15_45  = SHARE(GND)

	.dataa(!din_a[188]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_64 ),
	.sharein(Xd_0__inst_mult_12_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_43_sumout ),
	.cout(Xd_0__inst_mult_15_44 ),
	.shareout(Xd_0__inst_mult_15_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_93 (
// Equation(s):
// Xd_0__inst_mult_1_272  = SUM(( !Xd_0__inst_mult_1_392  $ (!Xd_0__inst_mult_1_396  $ (((din_b[16] & din_a[13])))) ) + ( Xd_0__inst_mult_1_258  ) + ( Xd_0__inst_mult_1_257  ))
// Xd_0__inst_mult_1_273  = CARRY(( !Xd_0__inst_mult_1_392  $ (!Xd_0__inst_mult_1_396  $ (((din_b[16] & din_a[13])))) ) + ( Xd_0__inst_mult_1_258  ) + ( Xd_0__inst_mult_1_257  ))
// Xd_0__inst_mult_1_274  = SHARE((!Xd_0__inst_mult_1_392  & (Xd_0__inst_mult_1_396  & (din_b[16] & din_a[13]))) # (Xd_0__inst_mult_1_392  & (((din_b[16] & din_a[13])) # (Xd_0__inst_mult_1_396 ))))

	.dataa(!Xd_0__inst_mult_1_392 ),
	.datab(!Xd_0__inst_mult_1_396 ),
	.datac(!din_b[16]),
	.datad(!din_a[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_257 ),
	.sharein(Xd_0__inst_mult_1_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_272 ),
	.cout(Xd_0__inst_mult_1_273 ),
	.shareout(Xd_0__inst_mult_1_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_94 (
// Equation(s):
// Xd_0__inst_mult_1_276  = SUM(( (din_a[12] & din_b[17]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_277  = CARRY(( (din_a[12] & din_b[17]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_278  = SHARE((din_a[12] & din_b[18]))

	.dataa(!din_a[12]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_276 ),
	.cout(Xd_0__inst_mult_1_277 ),
	.shareout(Xd_0__inst_mult_1_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_35 (
// Equation(s):
// Xd_0__inst_mult_0_35_sumout  = SUM(( (din_a[7] & din_b[0]) ) + ( Xd_0__inst_mult_1_65  ) + ( Xd_0__inst_mult_1_64  ))
// Xd_0__inst_mult_0_36  = CARRY(( (din_a[7] & din_b[0]) ) + ( Xd_0__inst_mult_1_65  ) + ( Xd_0__inst_mult_1_64  ))
// Xd_0__inst_mult_0_37  = SHARE(GND)

	.dataa(!din_a[7]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_64 ),
	.sharein(Xd_0__inst_mult_1_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_35_sumout ),
	.cout(Xd_0__inst_mult_0_36 ),
	.shareout(Xd_0__inst_mult_0_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_103 (
// Equation(s):
// Xd_0__inst_mult_12_324  = SUM(( !Xd_0__inst_mult_12_440  $ (!Xd_0__inst_mult_12_444 ) ) + ( Xd_0__inst_mult_12_318  ) + ( Xd_0__inst_mult_12_317  ))
// Xd_0__inst_mult_12_325  = CARRY(( !Xd_0__inst_mult_12_440  $ (!Xd_0__inst_mult_12_444 ) ) + ( Xd_0__inst_mult_12_318  ) + ( Xd_0__inst_mult_12_317  ))
// Xd_0__inst_mult_12_326  = SHARE((Xd_0__inst_mult_12_440  & Xd_0__inst_mult_12_444 ))

	.dataa(!Xd_0__inst_mult_12_440 ),
	.datab(!Xd_0__inst_mult_12_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_317 ),
	.sharein(Xd_0__inst_mult_12_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_324 ),
	.cout(Xd_0__inst_mult_12_325 ),
	.shareout(Xd_0__inst_mult_12_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_104 (
// Equation(s):
// Xd_0__inst_mult_12_328  = SUM(( (din_a[145] & din_b[149]) ) + ( Xd_0__inst_mult_12_322  ) + ( Xd_0__inst_mult_12_321  ))
// Xd_0__inst_mult_12_329  = CARRY(( (din_a[145] & din_b[149]) ) + ( Xd_0__inst_mult_12_322  ) + ( Xd_0__inst_mult_12_321  ))
// Xd_0__inst_mult_12_330  = SHARE((din_a[144] & din_b[151]))

	.dataa(!din_a[145]),
	.datab(!din_b[149]),
	.datac(!din_a[144]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_321 ),
	.sharein(Xd_0__inst_mult_12_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_328 ),
	.cout(Xd_0__inst_mult_12_329 ),
	.shareout(Xd_0__inst_mult_12_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_101 (
// Equation(s):
// Xd_0__inst_mult_13_304  = SUM(( !Xd_0__inst_mult_13_416  $ (!Xd_0__inst_mult_13_420 ) ) + ( Xd_0__inst_mult_13_298  ) + ( Xd_0__inst_mult_13_297  ))
// Xd_0__inst_mult_13_305  = CARRY(( !Xd_0__inst_mult_13_416  $ (!Xd_0__inst_mult_13_420 ) ) + ( Xd_0__inst_mult_13_298  ) + ( Xd_0__inst_mult_13_297  ))
// Xd_0__inst_mult_13_306  = SHARE((Xd_0__inst_mult_13_416  & Xd_0__inst_mult_13_420 ))

	.dataa(!Xd_0__inst_mult_13_416 ),
	.datab(!Xd_0__inst_mult_13_420 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_297 ),
	.sharein(Xd_0__inst_mult_13_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_304 ),
	.cout(Xd_0__inst_mult_13_305 ),
	.shareout(Xd_0__inst_mult_13_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_102 (
// Equation(s):
// Xd_0__inst_mult_13_308  = SUM(( (din_a[157] & din_b[161]) ) + ( Xd_0__inst_mult_13_302  ) + ( Xd_0__inst_mult_13_301  ))
// Xd_0__inst_mult_13_309  = CARRY(( (din_a[157] & din_b[161]) ) + ( Xd_0__inst_mult_13_302  ) + ( Xd_0__inst_mult_13_301  ))
// Xd_0__inst_mult_13_310  = SHARE((din_a[156] & din_b[163]))

	.dataa(!din_a[157]),
	.datab(!din_b[161]),
	.datac(!din_a[156]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_301 ),
	.sharein(Xd_0__inst_mult_13_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_308 ),
	.cout(Xd_0__inst_mult_13_309 ),
	.shareout(Xd_0__inst_mult_13_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_107 (
// Equation(s):
// Xd_0__inst_mult_14_328  = SUM(( !Xd_0__inst_mult_14_432  $ (!Xd_0__inst_mult_14_436 ) ) + ( Xd_0__inst_mult_14_322  ) + ( Xd_0__inst_mult_14_321  ))
// Xd_0__inst_mult_14_329  = CARRY(( !Xd_0__inst_mult_14_432  $ (!Xd_0__inst_mult_14_436 ) ) + ( Xd_0__inst_mult_14_322  ) + ( Xd_0__inst_mult_14_321  ))
// Xd_0__inst_mult_14_330  = SHARE((Xd_0__inst_mult_14_432  & Xd_0__inst_mult_14_436 ))

	.dataa(!Xd_0__inst_mult_14_432 ),
	.datab(!Xd_0__inst_mult_14_436 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_321 ),
	.sharein(Xd_0__inst_mult_14_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_328 ),
	.cout(Xd_0__inst_mult_14_329 ),
	.shareout(Xd_0__inst_mult_14_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_108 (
// Equation(s):
// Xd_0__inst_mult_14_332  = SUM(( (din_a[169] & din_b[173]) ) + ( Xd_0__inst_mult_14_326  ) + ( Xd_0__inst_mult_14_325  ))
// Xd_0__inst_mult_14_333  = CARRY(( (din_a[169] & din_b[173]) ) + ( Xd_0__inst_mult_14_326  ) + ( Xd_0__inst_mult_14_325  ))
// Xd_0__inst_mult_14_334  = SHARE((din_a[168] & din_b[175]))

	.dataa(!din_a[169]),
	.datab(!din_b[173]),
	.datac(!din_a[168]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_325 ),
	.sharein(Xd_0__inst_mult_14_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_332 ),
	.cout(Xd_0__inst_mult_14_333 ),
	.shareout(Xd_0__inst_mult_14_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_107 (
// Equation(s):
// Xd_0__inst_mult_15_328  = SUM(( !Xd_0__inst_mult_15_444  $ (!Xd_0__inst_mult_15_448 ) ) + ( Xd_0__inst_mult_15_322  ) + ( Xd_0__inst_mult_15_321  ))
// Xd_0__inst_mult_15_329  = CARRY(( !Xd_0__inst_mult_15_444  $ (!Xd_0__inst_mult_15_448 ) ) + ( Xd_0__inst_mult_15_322  ) + ( Xd_0__inst_mult_15_321  ))
// Xd_0__inst_mult_15_330  = SHARE((Xd_0__inst_mult_15_444  & Xd_0__inst_mult_15_448 ))

	.dataa(!Xd_0__inst_mult_15_444 ),
	.datab(!Xd_0__inst_mult_15_448 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_321 ),
	.sharein(Xd_0__inst_mult_15_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_328 ),
	.cout(Xd_0__inst_mult_15_329 ),
	.shareout(Xd_0__inst_mult_15_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_108 (
// Equation(s):
// Xd_0__inst_mult_15_332  = SUM(( (din_a[181] & din_b[185]) ) + ( Xd_0__inst_mult_15_326  ) + ( Xd_0__inst_mult_15_325  ))
// Xd_0__inst_mult_15_333  = CARRY(( (din_a[181] & din_b[185]) ) + ( Xd_0__inst_mult_15_326  ) + ( Xd_0__inst_mult_15_325  ))
// Xd_0__inst_mult_15_334  = SHARE((din_a[180] & din_b[187]))

	.dataa(!din_a[181]),
	.datab(!din_b[185]),
	.datac(!din_a[180]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_325 ),
	.sharein(Xd_0__inst_mult_15_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_332 ),
	.cout(Xd_0__inst_mult_15_333 ),
	.shareout(Xd_0__inst_mult_15_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_97 (
// Equation(s):
// Xd_0__inst_mult_10_300  = SUM(( !Xd_0__inst_mult_10_412  $ (!Xd_0__inst_mult_10_416 ) ) + ( Xd_0__inst_mult_10_294  ) + ( Xd_0__inst_mult_10_293  ))
// Xd_0__inst_mult_10_301  = CARRY(( !Xd_0__inst_mult_10_412  $ (!Xd_0__inst_mult_10_416 ) ) + ( Xd_0__inst_mult_10_294  ) + ( Xd_0__inst_mult_10_293  ))
// Xd_0__inst_mult_10_302  = SHARE((Xd_0__inst_mult_10_412  & Xd_0__inst_mult_10_416 ))

	.dataa(!Xd_0__inst_mult_10_412 ),
	.datab(!Xd_0__inst_mult_10_416 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_293 ),
	.sharein(Xd_0__inst_mult_10_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_300 ),
	.cout(Xd_0__inst_mult_10_301 ),
	.shareout(Xd_0__inst_mult_10_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_98 (
// Equation(s):
// Xd_0__inst_mult_10_304  = SUM(( (din_a[121] & din_b[125]) ) + ( Xd_0__inst_mult_10_298  ) + ( Xd_0__inst_mult_10_297  ))
// Xd_0__inst_mult_10_305  = CARRY(( (din_a[121] & din_b[125]) ) + ( Xd_0__inst_mult_10_298  ) + ( Xd_0__inst_mult_10_297  ))
// Xd_0__inst_mult_10_306  = SHARE((din_a[120] & din_b[127]))

	.dataa(!din_a[121]),
	.datab(!din_b[125]),
	.datac(!din_a[120]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_297 ),
	.sharein(Xd_0__inst_mult_10_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_304 ),
	.cout(Xd_0__inst_mult_10_305 ),
	.shareout(Xd_0__inst_mult_10_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_101 (
// Equation(s):
// Xd_0__inst_mult_11_304  = SUM(( !Xd_0__inst_mult_11_416  $ (!Xd_0__inst_mult_11_420 ) ) + ( Xd_0__inst_mult_11_298  ) + ( Xd_0__inst_mult_11_297  ))
// Xd_0__inst_mult_11_305  = CARRY(( !Xd_0__inst_mult_11_416  $ (!Xd_0__inst_mult_11_420 ) ) + ( Xd_0__inst_mult_11_298  ) + ( Xd_0__inst_mult_11_297  ))
// Xd_0__inst_mult_11_306  = SHARE((Xd_0__inst_mult_11_416  & Xd_0__inst_mult_11_420 ))

	.dataa(!Xd_0__inst_mult_11_416 ),
	.datab(!Xd_0__inst_mult_11_420 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_297 ),
	.sharein(Xd_0__inst_mult_11_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_304 ),
	.cout(Xd_0__inst_mult_11_305 ),
	.shareout(Xd_0__inst_mult_11_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_102 (
// Equation(s):
// Xd_0__inst_mult_11_308  = SUM(( (din_a[133] & din_b[137]) ) + ( Xd_0__inst_mult_11_302  ) + ( Xd_0__inst_mult_11_301  ))
// Xd_0__inst_mult_11_309  = CARRY(( (din_a[133] & din_b[137]) ) + ( Xd_0__inst_mult_11_302  ) + ( Xd_0__inst_mult_11_301  ))
// Xd_0__inst_mult_11_310  = SHARE((din_a[132] & din_b[139]))

	.dataa(!din_a[133]),
	.datab(!din_b[137]),
	.datac(!din_a[132]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_301 ),
	.sharein(Xd_0__inst_mult_11_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_308 ),
	.cout(Xd_0__inst_mult_11_309 ),
	.shareout(Xd_0__inst_mult_11_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_101 (
// Equation(s):
// Xd_0__inst_mult_8_304  = SUM(( !Xd_0__inst_mult_8_416  $ (!Xd_0__inst_mult_8_420 ) ) + ( Xd_0__inst_mult_8_298  ) + ( Xd_0__inst_mult_8_297  ))
// Xd_0__inst_mult_8_305  = CARRY(( !Xd_0__inst_mult_8_416  $ (!Xd_0__inst_mult_8_420 ) ) + ( Xd_0__inst_mult_8_298  ) + ( Xd_0__inst_mult_8_297  ))
// Xd_0__inst_mult_8_306  = SHARE((Xd_0__inst_mult_8_416  & Xd_0__inst_mult_8_420 ))

	.dataa(!Xd_0__inst_mult_8_416 ),
	.datab(!Xd_0__inst_mult_8_420 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_297 ),
	.sharein(Xd_0__inst_mult_8_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_304 ),
	.cout(Xd_0__inst_mult_8_305 ),
	.shareout(Xd_0__inst_mult_8_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_102 (
// Equation(s):
// Xd_0__inst_mult_8_308  = SUM(( (din_a[97] & din_b[101]) ) + ( Xd_0__inst_mult_8_302  ) + ( Xd_0__inst_mult_8_301  ))
// Xd_0__inst_mult_8_309  = CARRY(( (din_a[97] & din_b[101]) ) + ( Xd_0__inst_mult_8_302  ) + ( Xd_0__inst_mult_8_301  ))
// Xd_0__inst_mult_8_310  = SHARE((din_a[96] & din_b[103]))

	.dataa(!din_a[97]),
	.datab(!din_b[101]),
	.datac(!din_a[96]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_301 ),
	.sharein(Xd_0__inst_mult_8_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_308 ),
	.cout(Xd_0__inst_mult_8_309 ),
	.shareout(Xd_0__inst_mult_8_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_97 (
// Equation(s):
// Xd_0__inst_mult_9_300  = SUM(( !Xd_0__inst_mult_9_412  $ (!Xd_0__inst_mult_9_416 ) ) + ( Xd_0__inst_mult_9_294  ) + ( Xd_0__inst_mult_9_293  ))
// Xd_0__inst_mult_9_301  = CARRY(( !Xd_0__inst_mult_9_412  $ (!Xd_0__inst_mult_9_416 ) ) + ( Xd_0__inst_mult_9_294  ) + ( Xd_0__inst_mult_9_293  ))
// Xd_0__inst_mult_9_302  = SHARE((Xd_0__inst_mult_9_412  & Xd_0__inst_mult_9_416 ))

	.dataa(!Xd_0__inst_mult_9_412 ),
	.datab(!Xd_0__inst_mult_9_416 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_293 ),
	.sharein(Xd_0__inst_mult_9_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_300 ),
	.cout(Xd_0__inst_mult_9_301 ),
	.shareout(Xd_0__inst_mult_9_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_98 (
// Equation(s):
// Xd_0__inst_mult_9_304  = SUM(( (din_a[109] & din_b[113]) ) + ( Xd_0__inst_mult_9_298  ) + ( Xd_0__inst_mult_9_297  ))
// Xd_0__inst_mult_9_305  = CARRY(( (din_a[109] & din_b[113]) ) + ( Xd_0__inst_mult_9_298  ) + ( Xd_0__inst_mult_9_297  ))
// Xd_0__inst_mult_9_306  = SHARE((din_a[108] & din_b[115]))

	.dataa(!din_a[109]),
	.datab(!din_b[113]),
	.datac(!din_a[108]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_297 ),
	.sharein(Xd_0__inst_mult_9_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_304 ),
	.cout(Xd_0__inst_mult_9_305 ),
	.shareout(Xd_0__inst_mult_9_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_97 (
// Equation(s):
// Xd_0__inst_mult_6_300  = SUM(( !Xd_0__inst_mult_6_412  $ (!Xd_0__inst_mult_6_416 ) ) + ( Xd_0__inst_mult_6_294  ) + ( Xd_0__inst_mult_6_293  ))
// Xd_0__inst_mult_6_301  = CARRY(( !Xd_0__inst_mult_6_412  $ (!Xd_0__inst_mult_6_416 ) ) + ( Xd_0__inst_mult_6_294  ) + ( Xd_0__inst_mult_6_293  ))
// Xd_0__inst_mult_6_302  = SHARE((Xd_0__inst_mult_6_412  & Xd_0__inst_mult_6_416 ))

	.dataa(!Xd_0__inst_mult_6_412 ),
	.datab(!Xd_0__inst_mult_6_416 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_293 ),
	.sharein(Xd_0__inst_mult_6_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_300 ),
	.cout(Xd_0__inst_mult_6_301 ),
	.shareout(Xd_0__inst_mult_6_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_98 (
// Equation(s):
// Xd_0__inst_mult_6_304  = SUM(( (din_a[73] & din_b[77]) ) + ( Xd_0__inst_mult_6_298  ) + ( Xd_0__inst_mult_6_297  ))
// Xd_0__inst_mult_6_305  = CARRY(( (din_a[73] & din_b[77]) ) + ( Xd_0__inst_mult_6_298  ) + ( Xd_0__inst_mult_6_297  ))
// Xd_0__inst_mult_6_306  = SHARE((din_a[72] & din_b[79]))

	.dataa(!din_a[73]),
	.datab(!din_b[77]),
	.datac(!din_a[72]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_297 ),
	.sharein(Xd_0__inst_mult_6_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_304 ),
	.cout(Xd_0__inst_mult_6_305 ),
	.shareout(Xd_0__inst_mult_6_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_91 (
// Equation(s):
// Xd_0__inst_mult_7_276  = SUM(( !Xd_0__inst_mult_7_396  $ (!Xd_0__inst_mult_7_400 ) ) + ( Xd_0__inst_mult_7_270  ) + ( Xd_0__inst_mult_7_269  ))
// Xd_0__inst_mult_7_277  = CARRY(( !Xd_0__inst_mult_7_396  $ (!Xd_0__inst_mult_7_400 ) ) + ( Xd_0__inst_mult_7_270  ) + ( Xd_0__inst_mult_7_269  ))
// Xd_0__inst_mult_7_278  = SHARE((Xd_0__inst_mult_7_396  & Xd_0__inst_mult_7_400 ))

	.dataa(!Xd_0__inst_mult_7_396 ),
	.datab(!Xd_0__inst_mult_7_400 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_269 ),
	.sharein(Xd_0__inst_mult_7_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_276 ),
	.cout(Xd_0__inst_mult_7_277 ),
	.shareout(Xd_0__inst_mult_7_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_92 (
// Equation(s):
// Xd_0__inst_mult_7_280  = SUM(( (din_a[85] & din_b[89]) ) + ( Xd_0__inst_mult_7_274  ) + ( Xd_0__inst_mult_7_273  ))
// Xd_0__inst_mult_7_281  = CARRY(( (din_a[85] & din_b[89]) ) + ( Xd_0__inst_mult_7_274  ) + ( Xd_0__inst_mult_7_273  ))
// Xd_0__inst_mult_7_282  = SHARE((din_a[84] & din_b[91]))

	.dataa(!din_a[85]),
	.datab(!din_b[89]),
	.datac(!din_a[84]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_273 ),
	.sharein(Xd_0__inst_mult_7_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_280 ),
	.cout(Xd_0__inst_mult_7_281 ),
	.shareout(Xd_0__inst_mult_7_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_103 (
// Equation(s):
// Xd_0__inst_mult_4_312  = SUM(( !Xd_0__inst_mult_4_436  $ (!Xd_0__inst_mult_4_440 ) ) + ( Xd_0__inst_mult_4_306  ) + ( Xd_0__inst_mult_4_305  ))
// Xd_0__inst_mult_4_313  = CARRY(( !Xd_0__inst_mult_4_436  $ (!Xd_0__inst_mult_4_440 ) ) + ( Xd_0__inst_mult_4_306  ) + ( Xd_0__inst_mult_4_305  ))
// Xd_0__inst_mult_4_314  = SHARE((Xd_0__inst_mult_4_436  & Xd_0__inst_mult_4_440 ))

	.dataa(!Xd_0__inst_mult_4_436 ),
	.datab(!Xd_0__inst_mult_4_440 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_305 ),
	.sharein(Xd_0__inst_mult_4_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_312 ),
	.cout(Xd_0__inst_mult_4_313 ),
	.shareout(Xd_0__inst_mult_4_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_104 (
// Equation(s):
// Xd_0__inst_mult_4_316  = SUM(( (din_a[49] & din_b[53]) ) + ( Xd_0__inst_mult_4_310  ) + ( Xd_0__inst_mult_4_309  ))
// Xd_0__inst_mult_4_317  = CARRY(( (din_a[49] & din_b[53]) ) + ( Xd_0__inst_mult_4_310  ) + ( Xd_0__inst_mult_4_309  ))
// Xd_0__inst_mult_4_318  = SHARE((din_a[48] & din_b[55]))

	.dataa(!din_a[49]),
	.datab(!din_b[53]),
	.datac(!din_a[48]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_309 ),
	.sharein(Xd_0__inst_mult_4_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_316 ),
	.cout(Xd_0__inst_mult_4_317 ),
	.shareout(Xd_0__inst_mult_4_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_91 (
// Equation(s):
// Xd_0__inst_mult_5_276  = SUM(( !Xd_0__inst_mult_5_396  $ (!Xd_0__inst_mult_5_400 ) ) + ( Xd_0__inst_mult_5_270  ) + ( Xd_0__inst_mult_5_269  ))
// Xd_0__inst_mult_5_277  = CARRY(( !Xd_0__inst_mult_5_396  $ (!Xd_0__inst_mult_5_400 ) ) + ( Xd_0__inst_mult_5_270  ) + ( Xd_0__inst_mult_5_269  ))
// Xd_0__inst_mult_5_278  = SHARE((Xd_0__inst_mult_5_396  & Xd_0__inst_mult_5_400 ))

	.dataa(!Xd_0__inst_mult_5_396 ),
	.datab(!Xd_0__inst_mult_5_400 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_269 ),
	.sharein(Xd_0__inst_mult_5_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_276 ),
	.cout(Xd_0__inst_mult_5_277 ),
	.shareout(Xd_0__inst_mult_5_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_92 (
// Equation(s):
// Xd_0__inst_mult_5_280  = SUM(( (din_a[61] & din_b[65]) ) + ( Xd_0__inst_mult_5_274  ) + ( Xd_0__inst_mult_5_273  ))
// Xd_0__inst_mult_5_281  = CARRY(( (din_a[61] & din_b[65]) ) + ( Xd_0__inst_mult_5_274  ) + ( Xd_0__inst_mult_5_273  ))
// Xd_0__inst_mult_5_282  = SHARE((din_a[60] & din_b[67]))

	.dataa(!din_a[61]),
	.datab(!din_b[65]),
	.datac(!din_a[60]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_273 ),
	.sharein(Xd_0__inst_mult_5_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_280 ),
	.cout(Xd_0__inst_mult_5_281 ),
	.shareout(Xd_0__inst_mult_5_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_95 (
// Equation(s):
// Xd_0__inst_mult_2_280  = SUM(( !Xd_0__inst_mult_2_400  $ (!Xd_0__inst_mult_2_404 ) ) + ( Xd_0__inst_mult_2_274  ) + ( Xd_0__inst_mult_2_273  ))
// Xd_0__inst_mult_2_281  = CARRY(( !Xd_0__inst_mult_2_400  $ (!Xd_0__inst_mult_2_404 ) ) + ( Xd_0__inst_mult_2_274  ) + ( Xd_0__inst_mult_2_273  ))
// Xd_0__inst_mult_2_282  = SHARE((Xd_0__inst_mult_2_400  & Xd_0__inst_mult_2_404 ))

	.dataa(!Xd_0__inst_mult_2_400 ),
	.datab(!Xd_0__inst_mult_2_404 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_273 ),
	.sharein(Xd_0__inst_mult_2_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_280 ),
	.cout(Xd_0__inst_mult_2_281 ),
	.shareout(Xd_0__inst_mult_2_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_96 (
// Equation(s):
// Xd_0__inst_mult_2_284  = SUM(( (din_a[25] & din_b[29]) ) + ( Xd_0__inst_mult_2_278  ) + ( Xd_0__inst_mult_2_277  ))
// Xd_0__inst_mult_2_285  = CARRY(( (din_a[25] & din_b[29]) ) + ( Xd_0__inst_mult_2_278  ) + ( Xd_0__inst_mult_2_277  ))
// Xd_0__inst_mult_2_286  = SHARE((din_a[24] & din_b[31]))

	.dataa(!din_a[25]),
	.datab(!din_b[29]),
	.datac(!din_a[24]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_277 ),
	.sharein(Xd_0__inst_mult_2_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_284 ),
	.cout(Xd_0__inst_mult_2_285 ),
	.shareout(Xd_0__inst_mult_2_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_91 (
// Equation(s):
// Xd_0__inst_mult_3_276  = SUM(( !Xd_0__inst_mult_3_396  $ (!Xd_0__inst_mult_3_400 ) ) + ( Xd_0__inst_mult_3_270  ) + ( Xd_0__inst_mult_3_269  ))
// Xd_0__inst_mult_3_277  = CARRY(( !Xd_0__inst_mult_3_396  $ (!Xd_0__inst_mult_3_400 ) ) + ( Xd_0__inst_mult_3_270  ) + ( Xd_0__inst_mult_3_269  ))
// Xd_0__inst_mult_3_278  = SHARE((Xd_0__inst_mult_3_396  & Xd_0__inst_mult_3_400 ))

	.dataa(!Xd_0__inst_mult_3_396 ),
	.datab(!Xd_0__inst_mult_3_400 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_269 ),
	.sharein(Xd_0__inst_mult_3_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_276 ),
	.cout(Xd_0__inst_mult_3_277 ),
	.shareout(Xd_0__inst_mult_3_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_92 (
// Equation(s):
// Xd_0__inst_mult_3_280  = SUM(( (din_a[37] & din_b[41]) ) + ( Xd_0__inst_mult_3_274  ) + ( Xd_0__inst_mult_3_273  ))
// Xd_0__inst_mult_3_281  = CARRY(( (din_a[37] & din_b[41]) ) + ( Xd_0__inst_mult_3_274  ) + ( Xd_0__inst_mult_3_273  ))
// Xd_0__inst_mult_3_282  = SHARE((din_a[36] & din_b[43]))

	.dataa(!din_a[37]),
	.datab(!din_b[41]),
	.datac(!din_a[36]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_273 ),
	.sharein(Xd_0__inst_mult_3_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_280 ),
	.cout(Xd_0__inst_mult_3_281 ),
	.shareout(Xd_0__inst_mult_3_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_95 (
// Equation(s):
// Xd_0__inst_mult_0_280  = SUM(( !Xd_0__inst_mult_0_400  $ (!Xd_0__inst_mult_0_404 ) ) + ( Xd_0__inst_mult_0_274  ) + ( Xd_0__inst_mult_0_273  ))
// Xd_0__inst_mult_0_281  = CARRY(( !Xd_0__inst_mult_0_400  $ (!Xd_0__inst_mult_0_404 ) ) + ( Xd_0__inst_mult_0_274  ) + ( Xd_0__inst_mult_0_273  ))
// Xd_0__inst_mult_0_282  = SHARE((Xd_0__inst_mult_0_400  & Xd_0__inst_mult_0_404 ))

	.dataa(!Xd_0__inst_mult_0_400 ),
	.datab(!Xd_0__inst_mult_0_404 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_273 ),
	.sharein(Xd_0__inst_mult_0_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_280 ),
	.cout(Xd_0__inst_mult_0_281 ),
	.shareout(Xd_0__inst_mult_0_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_96 (
// Equation(s):
// Xd_0__inst_mult_0_284  = SUM(( (din_a[1] & din_b[5]) ) + ( Xd_0__inst_mult_0_278  ) + ( Xd_0__inst_mult_0_277  ))
// Xd_0__inst_mult_0_285  = CARRY(( (din_a[1] & din_b[5]) ) + ( Xd_0__inst_mult_0_278  ) + ( Xd_0__inst_mult_0_277  ))
// Xd_0__inst_mult_0_286  = SHARE((din_a[0] & din_b[7]))

	.dataa(!din_a[1]),
	.datab(!din_b[5]),
	.datac(!din_a[0]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_277 ),
	.sharein(Xd_0__inst_mult_0_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_284 ),
	.cout(Xd_0__inst_mult_0_285 ),
	.shareout(Xd_0__inst_mult_0_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_95 (
// Equation(s):
// Xd_0__inst_mult_1_280  = SUM(( !Xd_0__inst_mult_1_400  $ (!Xd_0__inst_mult_1_404 ) ) + ( Xd_0__inst_mult_1_274  ) + ( Xd_0__inst_mult_1_273  ))
// Xd_0__inst_mult_1_281  = CARRY(( !Xd_0__inst_mult_1_400  $ (!Xd_0__inst_mult_1_404 ) ) + ( Xd_0__inst_mult_1_274  ) + ( Xd_0__inst_mult_1_273  ))
// Xd_0__inst_mult_1_282  = SHARE((Xd_0__inst_mult_1_400  & Xd_0__inst_mult_1_404 ))

	.dataa(!Xd_0__inst_mult_1_400 ),
	.datab(!Xd_0__inst_mult_1_404 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_273 ),
	.sharein(Xd_0__inst_mult_1_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_280 ),
	.cout(Xd_0__inst_mult_1_281 ),
	.shareout(Xd_0__inst_mult_1_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_96 (
// Equation(s):
// Xd_0__inst_mult_1_284  = SUM(( (din_a[13] & din_b[17]) ) + ( Xd_0__inst_mult_1_278  ) + ( Xd_0__inst_mult_1_277  ))
// Xd_0__inst_mult_1_285  = CARRY(( (din_a[13] & din_b[17]) ) + ( Xd_0__inst_mult_1_278  ) + ( Xd_0__inst_mult_1_277  ))
// Xd_0__inst_mult_1_286  = SHARE((din_a[12] & din_b[19]))

	.dataa(!din_a[13]),
	.datab(!din_b[17]),
	.datac(!din_a[12]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_277 ),
	.sharein(Xd_0__inst_mult_1_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_284 ),
	.cout(Xd_0__inst_mult_1_285 ),
	.shareout(Xd_0__inst_mult_1_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_105 (
// Equation(s):
// Xd_0__inst_mult_12_332  = SUM(( !Xd_0__inst_mult_12_448  $ (!Xd_0__inst_mult_12_452  $ (Xd_0__inst_mult_12_43_sumout )) ) + ( Xd_0__inst_mult_12_326  ) + ( Xd_0__inst_mult_12_325  ))
// Xd_0__inst_mult_12_333  = CARRY(( !Xd_0__inst_mult_12_448  $ (!Xd_0__inst_mult_12_452  $ (Xd_0__inst_mult_12_43_sumout )) ) + ( Xd_0__inst_mult_12_326  ) + ( Xd_0__inst_mult_12_325  ))
// Xd_0__inst_mult_12_334  = SHARE((!Xd_0__inst_mult_12_448  & (Xd_0__inst_mult_12_452  & Xd_0__inst_mult_12_43_sumout )) # (Xd_0__inst_mult_12_448  & ((Xd_0__inst_mult_12_43_sumout ) # (Xd_0__inst_mult_12_452 ))))

	.dataa(!Xd_0__inst_mult_12_448 ),
	.datab(!Xd_0__inst_mult_12_452 ),
	.datac(!Xd_0__inst_mult_12_43_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_325 ),
	.sharein(Xd_0__inst_mult_12_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_332 ),
	.cout(Xd_0__inst_mult_12_333 ),
	.shareout(Xd_0__inst_mult_12_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_106 (
// Equation(s):
// Xd_0__inst_mult_12_336  = SUM(( (!din_a[145] & (((din_a[146] & din_b[149])))) # (din_a[145] & (!din_b[150] $ (((!din_a[146]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_12_330  ) + ( Xd_0__inst_mult_12_329  ))
// Xd_0__inst_mult_12_337  = CARRY(( (!din_a[145] & (((din_a[146] & din_b[149])))) # (din_a[145] & (!din_b[150] $ (((!din_a[146]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_12_330  ) + ( Xd_0__inst_mult_12_329  ))
// Xd_0__inst_mult_12_338  = SHARE((din_a[145] & (din_b[150] & (din_a[146] & din_b[149]))))

	.dataa(!din_a[145]),
	.datab(!din_b[150]),
	.datac(!din_a[146]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_329 ),
	.sharein(Xd_0__inst_mult_12_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_336 ),
	.cout(Xd_0__inst_mult_12_337 ),
	.shareout(Xd_0__inst_mult_12_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_103 (
// Equation(s):
// Xd_0__inst_mult_13_312  = SUM(( !Xd_0__inst_mult_13_424  $ (!Xd_0__inst_mult_13_428  $ (Xd_0__inst_mult_13_63_sumout )) ) + ( Xd_0__inst_mult_13_306  ) + ( Xd_0__inst_mult_13_305  ))
// Xd_0__inst_mult_13_313  = CARRY(( !Xd_0__inst_mult_13_424  $ (!Xd_0__inst_mult_13_428  $ (Xd_0__inst_mult_13_63_sumout )) ) + ( Xd_0__inst_mult_13_306  ) + ( Xd_0__inst_mult_13_305  ))
// Xd_0__inst_mult_13_314  = SHARE((!Xd_0__inst_mult_13_424  & (Xd_0__inst_mult_13_428  & Xd_0__inst_mult_13_63_sumout )) # (Xd_0__inst_mult_13_424  & ((Xd_0__inst_mult_13_63_sumout ) # (Xd_0__inst_mult_13_428 ))))

	.dataa(!Xd_0__inst_mult_13_424 ),
	.datab(!Xd_0__inst_mult_13_428 ),
	.datac(!Xd_0__inst_mult_13_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_305 ),
	.sharein(Xd_0__inst_mult_13_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_312 ),
	.cout(Xd_0__inst_mult_13_313 ),
	.shareout(Xd_0__inst_mult_13_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_104 (
// Equation(s):
// Xd_0__inst_mult_13_316  = SUM(( (!din_a[157] & (((din_a[158] & din_b[161])))) # (din_a[157] & (!din_b[162] $ (((!din_a[158]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_13_310  ) + ( Xd_0__inst_mult_13_309  ))
// Xd_0__inst_mult_13_317  = CARRY(( (!din_a[157] & (((din_a[158] & din_b[161])))) # (din_a[157] & (!din_b[162] $ (((!din_a[158]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_13_310  ) + ( Xd_0__inst_mult_13_309  ))
// Xd_0__inst_mult_13_318  = SHARE((din_a[157] & (din_b[162] & (din_a[158] & din_b[161]))))

	.dataa(!din_a[157]),
	.datab(!din_b[162]),
	.datac(!din_a[158]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_309 ),
	.sharein(Xd_0__inst_mult_13_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_316 ),
	.cout(Xd_0__inst_mult_13_317 ),
	.shareout(Xd_0__inst_mult_13_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_109 (
// Equation(s):
// Xd_0__inst_mult_14_336  = SUM(( !Xd_0__inst_mult_14_440  $ (!Xd_0__inst_mult_14_444  $ (Xd_0__inst_mult_14_35_sumout )) ) + ( Xd_0__inst_mult_14_330  ) + ( Xd_0__inst_mult_14_329  ))
// Xd_0__inst_mult_14_337  = CARRY(( !Xd_0__inst_mult_14_440  $ (!Xd_0__inst_mult_14_444  $ (Xd_0__inst_mult_14_35_sumout )) ) + ( Xd_0__inst_mult_14_330  ) + ( Xd_0__inst_mult_14_329  ))
// Xd_0__inst_mult_14_338  = SHARE((!Xd_0__inst_mult_14_440  & (Xd_0__inst_mult_14_444  & Xd_0__inst_mult_14_35_sumout )) # (Xd_0__inst_mult_14_440  & ((Xd_0__inst_mult_14_35_sumout ) # (Xd_0__inst_mult_14_444 ))))

	.dataa(!Xd_0__inst_mult_14_440 ),
	.datab(!Xd_0__inst_mult_14_444 ),
	.datac(!Xd_0__inst_mult_14_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_329 ),
	.sharein(Xd_0__inst_mult_14_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_336 ),
	.cout(Xd_0__inst_mult_14_337 ),
	.shareout(Xd_0__inst_mult_14_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_110 (
// Equation(s):
// Xd_0__inst_mult_14_340  = SUM(( (!din_a[169] & (((din_a[170] & din_b[173])))) # (din_a[169] & (!din_b[174] $ (((!din_a[170]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_14_334  ) + ( Xd_0__inst_mult_14_333  ))
// Xd_0__inst_mult_14_341  = CARRY(( (!din_a[169] & (((din_a[170] & din_b[173])))) # (din_a[169] & (!din_b[174] $ (((!din_a[170]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_14_334  ) + ( Xd_0__inst_mult_14_333  ))
// Xd_0__inst_mult_14_342  = SHARE((din_a[169] & (din_b[174] & (din_a[170] & din_b[173]))))

	.dataa(!din_a[169]),
	.datab(!din_b[174]),
	.datac(!din_a[170]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_333 ),
	.sharein(Xd_0__inst_mult_14_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_340 ),
	.cout(Xd_0__inst_mult_14_341 ),
	.shareout(Xd_0__inst_mult_14_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_109 (
// Equation(s):
// Xd_0__inst_mult_15_336  = SUM(( !Xd_0__inst_mult_15_452  $ (!Xd_0__inst_mult_15_456  $ (Xd_0__inst_mult_15_39_sumout )) ) + ( Xd_0__inst_mult_15_330  ) + ( Xd_0__inst_mult_15_329  ))
// Xd_0__inst_mult_15_337  = CARRY(( !Xd_0__inst_mult_15_452  $ (!Xd_0__inst_mult_15_456  $ (Xd_0__inst_mult_15_39_sumout )) ) + ( Xd_0__inst_mult_15_330  ) + ( Xd_0__inst_mult_15_329  ))
// Xd_0__inst_mult_15_338  = SHARE((!Xd_0__inst_mult_15_452  & (Xd_0__inst_mult_15_456  & Xd_0__inst_mult_15_39_sumout )) # (Xd_0__inst_mult_15_452  & ((Xd_0__inst_mult_15_39_sumout ) # (Xd_0__inst_mult_15_456 ))))

	.dataa(!Xd_0__inst_mult_15_452 ),
	.datab(!Xd_0__inst_mult_15_456 ),
	.datac(!Xd_0__inst_mult_15_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_329 ),
	.sharein(Xd_0__inst_mult_15_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_336 ),
	.cout(Xd_0__inst_mult_15_337 ),
	.shareout(Xd_0__inst_mult_15_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_110 (
// Equation(s):
// Xd_0__inst_mult_15_340  = SUM(( (!din_a[181] & (((din_a[182] & din_b[185])))) # (din_a[181] & (!din_b[186] $ (((!din_a[182]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_15_334  ) + ( Xd_0__inst_mult_15_333  ))
// Xd_0__inst_mult_15_341  = CARRY(( (!din_a[181] & (((din_a[182] & din_b[185])))) # (din_a[181] & (!din_b[186] $ (((!din_a[182]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_15_334  ) + ( Xd_0__inst_mult_15_333  ))
// Xd_0__inst_mult_15_342  = SHARE((din_a[181] & (din_b[186] & (din_a[182] & din_b[185]))))

	.dataa(!din_a[181]),
	.datab(!din_b[186]),
	.datac(!din_a[182]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_333 ),
	.sharein(Xd_0__inst_mult_15_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_340 ),
	.cout(Xd_0__inst_mult_15_341 ),
	.shareout(Xd_0__inst_mult_15_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_99 (
// Equation(s):
// Xd_0__inst_mult_10_308  = SUM(( !Xd_0__inst_mult_10_420  $ (!Xd_0__inst_mult_10_424  $ (Xd_0__inst_mult_10_35_sumout )) ) + ( Xd_0__inst_mult_10_302  ) + ( Xd_0__inst_mult_10_301  ))
// Xd_0__inst_mult_10_309  = CARRY(( !Xd_0__inst_mult_10_420  $ (!Xd_0__inst_mult_10_424  $ (Xd_0__inst_mult_10_35_sumout )) ) + ( Xd_0__inst_mult_10_302  ) + ( Xd_0__inst_mult_10_301  ))
// Xd_0__inst_mult_10_310  = SHARE((!Xd_0__inst_mult_10_420  & (Xd_0__inst_mult_10_424  & Xd_0__inst_mult_10_35_sumout )) # (Xd_0__inst_mult_10_420  & ((Xd_0__inst_mult_10_35_sumout ) # (Xd_0__inst_mult_10_424 ))))

	.dataa(!Xd_0__inst_mult_10_420 ),
	.datab(!Xd_0__inst_mult_10_424 ),
	.datac(!Xd_0__inst_mult_10_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_301 ),
	.sharein(Xd_0__inst_mult_10_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_308 ),
	.cout(Xd_0__inst_mult_10_309 ),
	.shareout(Xd_0__inst_mult_10_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_100 (
// Equation(s):
// Xd_0__inst_mult_10_312  = SUM(( (!din_a[121] & (((din_a[122] & din_b[125])))) # (din_a[121] & (!din_b[126] $ (((!din_a[122]) # (!din_b[125]))))) ) + ( Xd_0__inst_mult_10_306  ) + ( Xd_0__inst_mult_10_305  ))
// Xd_0__inst_mult_10_313  = CARRY(( (!din_a[121] & (((din_a[122] & din_b[125])))) # (din_a[121] & (!din_b[126] $ (((!din_a[122]) # (!din_b[125]))))) ) + ( Xd_0__inst_mult_10_306  ) + ( Xd_0__inst_mult_10_305  ))
// Xd_0__inst_mult_10_314  = SHARE((din_a[121] & (din_b[126] & (din_a[122] & din_b[125]))))

	.dataa(!din_a[121]),
	.datab(!din_b[126]),
	.datac(!din_a[122]),
	.datad(!din_b[125]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_305 ),
	.sharein(Xd_0__inst_mult_10_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_312 ),
	.cout(Xd_0__inst_mult_10_313 ),
	.shareout(Xd_0__inst_mult_10_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_103 (
// Equation(s):
// Xd_0__inst_mult_11_312  = SUM(( !Xd_0__inst_mult_11_424  $ (!Xd_0__inst_mult_11_428  $ (Xd_0__inst_mult_11_63_sumout )) ) + ( Xd_0__inst_mult_11_306  ) + ( Xd_0__inst_mult_11_305  ))
// Xd_0__inst_mult_11_313  = CARRY(( !Xd_0__inst_mult_11_424  $ (!Xd_0__inst_mult_11_428  $ (Xd_0__inst_mult_11_63_sumout )) ) + ( Xd_0__inst_mult_11_306  ) + ( Xd_0__inst_mult_11_305  ))
// Xd_0__inst_mult_11_314  = SHARE((!Xd_0__inst_mult_11_424  & (Xd_0__inst_mult_11_428  & Xd_0__inst_mult_11_63_sumout )) # (Xd_0__inst_mult_11_424  & ((Xd_0__inst_mult_11_63_sumout ) # (Xd_0__inst_mult_11_428 ))))

	.dataa(!Xd_0__inst_mult_11_424 ),
	.datab(!Xd_0__inst_mult_11_428 ),
	.datac(!Xd_0__inst_mult_11_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_305 ),
	.sharein(Xd_0__inst_mult_11_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_312 ),
	.cout(Xd_0__inst_mult_11_313 ),
	.shareout(Xd_0__inst_mult_11_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_104 (
// Equation(s):
// Xd_0__inst_mult_11_316  = SUM(( (!din_a[133] & (((din_a[134] & din_b[137])))) # (din_a[133] & (!din_b[138] $ (((!din_a[134]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_11_310  ) + ( Xd_0__inst_mult_11_309  ))
// Xd_0__inst_mult_11_317  = CARRY(( (!din_a[133] & (((din_a[134] & din_b[137])))) # (din_a[133] & (!din_b[138] $ (((!din_a[134]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_11_310  ) + ( Xd_0__inst_mult_11_309  ))
// Xd_0__inst_mult_11_318  = SHARE((din_a[133] & (din_b[138] & (din_a[134] & din_b[137]))))

	.dataa(!din_a[133]),
	.datab(!din_b[138]),
	.datac(!din_a[134]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_309 ),
	.sharein(Xd_0__inst_mult_11_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_316 ),
	.cout(Xd_0__inst_mult_11_317 ),
	.shareout(Xd_0__inst_mult_11_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_103 (
// Equation(s):
// Xd_0__inst_mult_8_312  = SUM(( !Xd_0__inst_mult_8_424  $ (!Xd_0__inst_mult_8_428  $ (Xd_0__inst_mult_8_63_sumout )) ) + ( Xd_0__inst_mult_8_306  ) + ( Xd_0__inst_mult_8_305  ))
// Xd_0__inst_mult_8_313  = CARRY(( !Xd_0__inst_mult_8_424  $ (!Xd_0__inst_mult_8_428  $ (Xd_0__inst_mult_8_63_sumout )) ) + ( Xd_0__inst_mult_8_306  ) + ( Xd_0__inst_mult_8_305  ))
// Xd_0__inst_mult_8_314  = SHARE((!Xd_0__inst_mult_8_424  & (Xd_0__inst_mult_8_428  & Xd_0__inst_mult_8_63_sumout )) # (Xd_0__inst_mult_8_424  & ((Xd_0__inst_mult_8_63_sumout ) # (Xd_0__inst_mult_8_428 ))))

	.dataa(!Xd_0__inst_mult_8_424 ),
	.datab(!Xd_0__inst_mult_8_428 ),
	.datac(!Xd_0__inst_mult_8_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_305 ),
	.sharein(Xd_0__inst_mult_8_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_312 ),
	.cout(Xd_0__inst_mult_8_313 ),
	.shareout(Xd_0__inst_mult_8_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_104 (
// Equation(s):
// Xd_0__inst_mult_8_316  = SUM(( (!din_a[97] & (((din_a[98] & din_b[101])))) # (din_a[97] & (!din_b[102] $ (((!din_a[98]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_8_310  ) + ( Xd_0__inst_mult_8_309  ))
// Xd_0__inst_mult_8_317  = CARRY(( (!din_a[97] & (((din_a[98] & din_b[101])))) # (din_a[97] & (!din_b[102] $ (((!din_a[98]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_8_310  ) + ( Xd_0__inst_mult_8_309  ))
// Xd_0__inst_mult_8_318  = SHARE((din_a[97] & (din_b[102] & (din_a[98] & din_b[101]))))

	.dataa(!din_a[97]),
	.datab(!din_b[102]),
	.datac(!din_a[98]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_309 ),
	.sharein(Xd_0__inst_mult_8_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_316 ),
	.cout(Xd_0__inst_mult_8_317 ),
	.shareout(Xd_0__inst_mult_8_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_99 (
// Equation(s):
// Xd_0__inst_mult_9_308  = SUM(( !Xd_0__inst_mult_9_420  $ (!Xd_0__inst_mult_9_424  $ (Xd_0__inst_mult_9_59_sumout )) ) + ( Xd_0__inst_mult_9_302  ) + ( Xd_0__inst_mult_9_301  ))
// Xd_0__inst_mult_9_309  = CARRY(( !Xd_0__inst_mult_9_420  $ (!Xd_0__inst_mult_9_424  $ (Xd_0__inst_mult_9_59_sumout )) ) + ( Xd_0__inst_mult_9_302  ) + ( Xd_0__inst_mult_9_301  ))
// Xd_0__inst_mult_9_310  = SHARE((!Xd_0__inst_mult_9_420  & (Xd_0__inst_mult_9_424  & Xd_0__inst_mult_9_59_sumout )) # (Xd_0__inst_mult_9_420  & ((Xd_0__inst_mult_9_59_sumout ) # (Xd_0__inst_mult_9_424 ))))

	.dataa(!Xd_0__inst_mult_9_420 ),
	.datab(!Xd_0__inst_mult_9_424 ),
	.datac(!Xd_0__inst_mult_9_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_301 ),
	.sharein(Xd_0__inst_mult_9_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_308 ),
	.cout(Xd_0__inst_mult_9_309 ),
	.shareout(Xd_0__inst_mult_9_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_100 (
// Equation(s):
// Xd_0__inst_mult_9_312  = SUM(( (!din_a[109] & (((din_a[110] & din_b[113])))) # (din_a[109] & (!din_b[114] $ (((!din_a[110]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_9_306  ) + ( Xd_0__inst_mult_9_305  ))
// Xd_0__inst_mult_9_313  = CARRY(( (!din_a[109] & (((din_a[110] & din_b[113])))) # (din_a[109] & (!din_b[114] $ (((!din_a[110]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_9_306  ) + ( Xd_0__inst_mult_9_305  ))
// Xd_0__inst_mult_9_314  = SHARE((din_a[109] & (din_b[114] & (din_a[110] & din_b[113]))))

	.dataa(!din_a[109]),
	.datab(!din_b[114]),
	.datac(!din_a[110]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_305 ),
	.sharein(Xd_0__inst_mult_9_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_312 ),
	.cout(Xd_0__inst_mult_9_313 ),
	.shareout(Xd_0__inst_mult_9_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_99 (
// Equation(s):
// Xd_0__inst_mult_6_308  = SUM(( !Xd_0__inst_mult_6_420  $ (!Xd_0__inst_mult_6_424  $ (Xd_0__inst_mult_6_59_sumout )) ) + ( Xd_0__inst_mult_6_302  ) + ( Xd_0__inst_mult_6_301  ))
// Xd_0__inst_mult_6_309  = CARRY(( !Xd_0__inst_mult_6_420  $ (!Xd_0__inst_mult_6_424  $ (Xd_0__inst_mult_6_59_sumout )) ) + ( Xd_0__inst_mult_6_302  ) + ( Xd_0__inst_mult_6_301  ))
// Xd_0__inst_mult_6_310  = SHARE((!Xd_0__inst_mult_6_420  & (Xd_0__inst_mult_6_424  & Xd_0__inst_mult_6_59_sumout )) # (Xd_0__inst_mult_6_420  & ((Xd_0__inst_mult_6_59_sumout ) # (Xd_0__inst_mult_6_424 ))))

	.dataa(!Xd_0__inst_mult_6_420 ),
	.datab(!Xd_0__inst_mult_6_424 ),
	.datac(!Xd_0__inst_mult_6_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_301 ),
	.sharein(Xd_0__inst_mult_6_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_308 ),
	.cout(Xd_0__inst_mult_6_309 ),
	.shareout(Xd_0__inst_mult_6_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_100 (
// Equation(s):
// Xd_0__inst_mult_6_312  = SUM(( (!din_a[73] & (((din_a[74] & din_b[77])))) # (din_a[73] & (!din_b[78] $ (((!din_a[74]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_306  ) + ( Xd_0__inst_mult_6_305  ))
// Xd_0__inst_mult_6_313  = CARRY(( (!din_a[73] & (((din_a[74] & din_b[77])))) # (din_a[73] & (!din_b[78] $ (((!din_a[74]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_306  ) + ( Xd_0__inst_mult_6_305  ))
// Xd_0__inst_mult_6_314  = SHARE((din_a[73] & (din_b[78] & (din_a[74] & din_b[77]))))

	.dataa(!din_a[73]),
	.datab(!din_b[78]),
	.datac(!din_a[74]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_305 ),
	.sharein(Xd_0__inst_mult_6_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_312 ),
	.cout(Xd_0__inst_mult_6_313 ),
	.shareout(Xd_0__inst_mult_6_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_93 (
// Equation(s):
// Xd_0__inst_mult_7_284  = SUM(( !Xd_0__inst_mult_7_404  $ (!Xd_0__inst_mult_7_408  $ (Xd_0__inst_mult_7_55_sumout )) ) + ( Xd_0__inst_mult_7_278  ) + ( Xd_0__inst_mult_7_277  ))
// Xd_0__inst_mult_7_285  = CARRY(( !Xd_0__inst_mult_7_404  $ (!Xd_0__inst_mult_7_408  $ (Xd_0__inst_mult_7_55_sumout )) ) + ( Xd_0__inst_mult_7_278  ) + ( Xd_0__inst_mult_7_277  ))
// Xd_0__inst_mult_7_286  = SHARE((!Xd_0__inst_mult_7_404  & (Xd_0__inst_mult_7_408  & Xd_0__inst_mult_7_55_sumout )) # (Xd_0__inst_mult_7_404  & ((Xd_0__inst_mult_7_55_sumout ) # (Xd_0__inst_mult_7_408 ))))

	.dataa(!Xd_0__inst_mult_7_404 ),
	.datab(!Xd_0__inst_mult_7_408 ),
	.datac(!Xd_0__inst_mult_7_55_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_277 ),
	.sharein(Xd_0__inst_mult_7_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_284 ),
	.cout(Xd_0__inst_mult_7_285 ),
	.shareout(Xd_0__inst_mult_7_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_94 (
// Equation(s):
// Xd_0__inst_mult_7_288  = SUM(( (!din_a[85] & (((din_a[86] & din_b[89])))) # (din_a[85] & (!din_b[90] $ (((!din_a[86]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_282  ) + ( Xd_0__inst_mult_7_281  ))
// Xd_0__inst_mult_7_289  = CARRY(( (!din_a[85] & (((din_a[86] & din_b[89])))) # (din_a[85] & (!din_b[90] $ (((!din_a[86]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_282  ) + ( Xd_0__inst_mult_7_281  ))
// Xd_0__inst_mult_7_290  = SHARE((din_a[85] & (din_b[90] & (din_a[86] & din_b[89]))))

	.dataa(!din_a[85]),
	.datab(!din_b[90]),
	.datac(!din_a[86]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_281 ),
	.sharein(Xd_0__inst_mult_7_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_288 ),
	.cout(Xd_0__inst_mult_7_289 ),
	.shareout(Xd_0__inst_mult_7_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_105 (
// Equation(s):
// Xd_0__inst_mult_4_320  = SUM(( !Xd_0__inst_mult_4_444  $ (!Xd_0__inst_mult_4_448  $ (Xd_0__inst_mult_4_59_sumout )) ) + ( Xd_0__inst_mult_4_314  ) + ( Xd_0__inst_mult_4_313  ))
// Xd_0__inst_mult_4_321  = CARRY(( !Xd_0__inst_mult_4_444  $ (!Xd_0__inst_mult_4_448  $ (Xd_0__inst_mult_4_59_sumout )) ) + ( Xd_0__inst_mult_4_314  ) + ( Xd_0__inst_mult_4_313  ))
// Xd_0__inst_mult_4_322  = SHARE((!Xd_0__inst_mult_4_444  & (Xd_0__inst_mult_4_448  & Xd_0__inst_mult_4_59_sumout )) # (Xd_0__inst_mult_4_444  & ((Xd_0__inst_mult_4_59_sumout ) # (Xd_0__inst_mult_4_448 ))))

	.dataa(!Xd_0__inst_mult_4_444 ),
	.datab(!Xd_0__inst_mult_4_448 ),
	.datac(!Xd_0__inst_mult_4_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_313 ),
	.sharein(Xd_0__inst_mult_4_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_320 ),
	.cout(Xd_0__inst_mult_4_321 ),
	.shareout(Xd_0__inst_mult_4_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_106 (
// Equation(s):
// Xd_0__inst_mult_4_324  = SUM(( (!din_a[49] & (((din_a[50] & din_b[53])))) # (din_a[49] & (!din_b[54] $ (((!din_a[50]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_318  ) + ( Xd_0__inst_mult_4_317  ))
// Xd_0__inst_mult_4_325  = CARRY(( (!din_a[49] & (((din_a[50] & din_b[53])))) # (din_a[49] & (!din_b[54] $ (((!din_a[50]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_318  ) + ( Xd_0__inst_mult_4_317  ))
// Xd_0__inst_mult_4_326  = SHARE((din_a[49] & (din_b[54] & (din_a[50] & din_b[53]))))

	.dataa(!din_a[49]),
	.datab(!din_b[54]),
	.datac(!din_a[50]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_317 ),
	.sharein(Xd_0__inst_mult_4_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_324 ),
	.cout(Xd_0__inst_mult_4_325 ),
	.shareout(Xd_0__inst_mult_4_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_93 (
// Equation(s):
// Xd_0__inst_mult_5_284  = SUM(( !Xd_0__inst_mult_5_404  $ (!Xd_0__inst_mult_5_408  $ (Xd_0__inst_mult_5_59_sumout )) ) + ( Xd_0__inst_mult_5_278  ) + ( Xd_0__inst_mult_5_277  ))
// Xd_0__inst_mult_5_285  = CARRY(( !Xd_0__inst_mult_5_404  $ (!Xd_0__inst_mult_5_408  $ (Xd_0__inst_mult_5_59_sumout )) ) + ( Xd_0__inst_mult_5_278  ) + ( Xd_0__inst_mult_5_277  ))
// Xd_0__inst_mult_5_286  = SHARE((!Xd_0__inst_mult_5_404  & (Xd_0__inst_mult_5_408  & Xd_0__inst_mult_5_59_sumout )) # (Xd_0__inst_mult_5_404  & ((Xd_0__inst_mult_5_59_sumout ) # (Xd_0__inst_mult_5_408 ))))

	.dataa(!Xd_0__inst_mult_5_404 ),
	.datab(!Xd_0__inst_mult_5_408 ),
	.datac(!Xd_0__inst_mult_5_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_277 ),
	.sharein(Xd_0__inst_mult_5_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_284 ),
	.cout(Xd_0__inst_mult_5_285 ),
	.shareout(Xd_0__inst_mult_5_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_94 (
// Equation(s):
// Xd_0__inst_mult_5_288  = SUM(( (!din_a[61] & (((din_a[62] & din_b[65])))) # (din_a[61] & (!din_b[66] $ (((!din_a[62]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_282  ) + ( Xd_0__inst_mult_5_281  ))
// Xd_0__inst_mult_5_289  = CARRY(( (!din_a[61] & (((din_a[62] & din_b[65])))) # (din_a[61] & (!din_b[66] $ (((!din_a[62]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_282  ) + ( Xd_0__inst_mult_5_281  ))
// Xd_0__inst_mult_5_290  = SHARE((din_a[61] & (din_b[66] & (din_a[62] & din_b[65]))))

	.dataa(!din_a[61]),
	.datab(!din_b[66]),
	.datac(!din_a[62]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_281 ),
	.sharein(Xd_0__inst_mult_5_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_288 ),
	.cout(Xd_0__inst_mult_5_289 ),
	.shareout(Xd_0__inst_mult_5_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_97 (
// Equation(s):
// Xd_0__inst_mult_2_288  = SUM(( !Xd_0__inst_mult_2_408  $ (!Xd_0__inst_mult_2_412  $ (Xd_0__inst_mult_2_59_sumout )) ) + ( Xd_0__inst_mult_2_282  ) + ( Xd_0__inst_mult_2_281  ))
// Xd_0__inst_mult_2_289  = CARRY(( !Xd_0__inst_mult_2_408  $ (!Xd_0__inst_mult_2_412  $ (Xd_0__inst_mult_2_59_sumout )) ) + ( Xd_0__inst_mult_2_282  ) + ( Xd_0__inst_mult_2_281  ))
// Xd_0__inst_mult_2_290  = SHARE((!Xd_0__inst_mult_2_408  & (Xd_0__inst_mult_2_412  & Xd_0__inst_mult_2_59_sumout )) # (Xd_0__inst_mult_2_408  & ((Xd_0__inst_mult_2_59_sumout ) # (Xd_0__inst_mult_2_412 ))))

	.dataa(!Xd_0__inst_mult_2_408 ),
	.datab(!Xd_0__inst_mult_2_412 ),
	.datac(!Xd_0__inst_mult_2_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_281 ),
	.sharein(Xd_0__inst_mult_2_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_288 ),
	.cout(Xd_0__inst_mult_2_289 ),
	.shareout(Xd_0__inst_mult_2_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_98 (
// Equation(s):
// Xd_0__inst_mult_2_292  = SUM(( (!din_a[25] & (((din_a[26] & din_b[29])))) # (din_a[25] & (!din_b[30] $ (((!din_a[26]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_286  ) + ( Xd_0__inst_mult_2_285  ))
// Xd_0__inst_mult_2_293  = CARRY(( (!din_a[25] & (((din_a[26] & din_b[29])))) # (din_a[25] & (!din_b[30] $ (((!din_a[26]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_286  ) + ( Xd_0__inst_mult_2_285  ))
// Xd_0__inst_mult_2_294  = SHARE((din_a[25] & (din_b[30] & (din_a[26] & din_b[29]))))

	.dataa(!din_a[25]),
	.datab(!din_b[30]),
	.datac(!din_a[26]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_285 ),
	.sharein(Xd_0__inst_mult_2_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_292 ),
	.cout(Xd_0__inst_mult_2_293 ),
	.shareout(Xd_0__inst_mult_2_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_93 (
// Equation(s):
// Xd_0__inst_mult_3_284  = SUM(( !Xd_0__inst_mult_3_404  $ (!Xd_0__inst_mult_3_408  $ (Xd_0__inst_mult_3_35_sumout )) ) + ( Xd_0__inst_mult_3_278  ) + ( Xd_0__inst_mult_3_277  ))
// Xd_0__inst_mult_3_285  = CARRY(( !Xd_0__inst_mult_3_404  $ (!Xd_0__inst_mult_3_408  $ (Xd_0__inst_mult_3_35_sumout )) ) + ( Xd_0__inst_mult_3_278  ) + ( Xd_0__inst_mult_3_277  ))
// Xd_0__inst_mult_3_286  = SHARE((!Xd_0__inst_mult_3_404  & (Xd_0__inst_mult_3_408  & Xd_0__inst_mult_3_35_sumout )) # (Xd_0__inst_mult_3_404  & ((Xd_0__inst_mult_3_35_sumout ) # (Xd_0__inst_mult_3_408 ))))

	.dataa(!Xd_0__inst_mult_3_404 ),
	.datab(!Xd_0__inst_mult_3_408 ),
	.datac(!Xd_0__inst_mult_3_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_277 ),
	.sharein(Xd_0__inst_mult_3_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_284 ),
	.cout(Xd_0__inst_mult_3_285 ),
	.shareout(Xd_0__inst_mult_3_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_94 (
// Equation(s):
// Xd_0__inst_mult_3_288  = SUM(( (!din_a[37] & (((din_a[38] & din_b[41])))) # (din_a[37] & (!din_b[42] $ (((!din_a[38]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_282  ) + ( Xd_0__inst_mult_3_281  ))
// Xd_0__inst_mult_3_289  = CARRY(( (!din_a[37] & (((din_a[38] & din_b[41])))) # (din_a[37] & (!din_b[42] $ (((!din_a[38]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_282  ) + ( Xd_0__inst_mult_3_281  ))
// Xd_0__inst_mult_3_290  = SHARE((din_a[37] & (din_b[42] & (din_a[38] & din_b[41]))))

	.dataa(!din_a[37]),
	.datab(!din_b[42]),
	.datac(!din_a[38]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_281 ),
	.sharein(Xd_0__inst_mult_3_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_288 ),
	.cout(Xd_0__inst_mult_3_289 ),
	.shareout(Xd_0__inst_mult_3_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_97 (
// Equation(s):
// Xd_0__inst_mult_0_288  = SUM(( !Xd_0__inst_mult_0_408  $ (!Xd_0__inst_mult_0_412  $ (Xd_0__inst_mult_0_35_sumout )) ) + ( Xd_0__inst_mult_0_282  ) + ( Xd_0__inst_mult_0_281  ))
// Xd_0__inst_mult_0_289  = CARRY(( !Xd_0__inst_mult_0_408  $ (!Xd_0__inst_mult_0_412  $ (Xd_0__inst_mult_0_35_sumout )) ) + ( Xd_0__inst_mult_0_282  ) + ( Xd_0__inst_mult_0_281  ))
// Xd_0__inst_mult_0_290  = SHARE((!Xd_0__inst_mult_0_408  & (Xd_0__inst_mult_0_412  & Xd_0__inst_mult_0_35_sumout )) # (Xd_0__inst_mult_0_408  & ((Xd_0__inst_mult_0_35_sumout ) # (Xd_0__inst_mult_0_412 ))))

	.dataa(!Xd_0__inst_mult_0_408 ),
	.datab(!Xd_0__inst_mult_0_412 ),
	.datac(!Xd_0__inst_mult_0_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_281 ),
	.sharein(Xd_0__inst_mult_0_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_288 ),
	.cout(Xd_0__inst_mult_0_289 ),
	.shareout(Xd_0__inst_mult_0_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_98 (
// Equation(s):
// Xd_0__inst_mult_0_292  = SUM(( (!din_a[1] & (((din_a[2] & din_b[5])))) # (din_a[1] & (!din_b[6] $ (((!din_a[2]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_286  ) + ( Xd_0__inst_mult_0_285  ))
// Xd_0__inst_mult_0_293  = CARRY(( (!din_a[1] & (((din_a[2] & din_b[5])))) # (din_a[1] & (!din_b[6] $ (((!din_a[2]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_286  ) + ( Xd_0__inst_mult_0_285  ))
// Xd_0__inst_mult_0_294  = SHARE((din_a[1] & (din_b[6] & (din_a[2] & din_b[5]))))

	.dataa(!din_a[1]),
	.datab(!din_b[6]),
	.datac(!din_a[2]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_285 ),
	.sharein(Xd_0__inst_mult_0_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_292 ),
	.cout(Xd_0__inst_mult_0_293 ),
	.shareout(Xd_0__inst_mult_0_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_97 (
// Equation(s):
// Xd_0__inst_mult_1_288  = SUM(( !Xd_0__inst_mult_1_408  $ (!Xd_0__inst_mult_1_412  $ (Xd_0__inst_mult_1_63_sumout )) ) + ( Xd_0__inst_mult_1_282  ) + ( Xd_0__inst_mult_1_281  ))
// Xd_0__inst_mult_1_289  = CARRY(( !Xd_0__inst_mult_1_408  $ (!Xd_0__inst_mult_1_412  $ (Xd_0__inst_mult_1_63_sumout )) ) + ( Xd_0__inst_mult_1_282  ) + ( Xd_0__inst_mult_1_281  ))
// Xd_0__inst_mult_1_290  = SHARE((!Xd_0__inst_mult_1_408  & (Xd_0__inst_mult_1_412  & Xd_0__inst_mult_1_63_sumout )) # (Xd_0__inst_mult_1_408  & ((Xd_0__inst_mult_1_63_sumout ) # (Xd_0__inst_mult_1_412 ))))

	.dataa(!Xd_0__inst_mult_1_408 ),
	.datab(!Xd_0__inst_mult_1_412 ),
	.datac(!Xd_0__inst_mult_1_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_281 ),
	.sharein(Xd_0__inst_mult_1_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_288 ),
	.cout(Xd_0__inst_mult_1_289 ),
	.shareout(Xd_0__inst_mult_1_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_98 (
// Equation(s):
// Xd_0__inst_mult_1_292  = SUM(( (!din_a[13] & (((din_a[14] & din_b[17])))) # (din_a[13] & (!din_b[18] $ (((!din_a[14]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_286  ) + ( Xd_0__inst_mult_1_285  ))
// Xd_0__inst_mult_1_293  = CARRY(( (!din_a[13] & (((din_a[14] & din_b[17])))) # (din_a[13] & (!din_b[18] $ (((!din_a[14]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_286  ) + ( Xd_0__inst_mult_1_285  ))
// Xd_0__inst_mult_1_294  = SHARE((din_a[13] & (din_b[18] & (din_a[14] & din_b[17]))))

	.dataa(!din_a[13]),
	.datab(!din_b[18]),
	.datac(!din_a[14]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_285 ),
	.sharein(Xd_0__inst_mult_1_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_292 ),
	.cout(Xd_0__inst_mult_1_293 ),
	.shareout(Xd_0__inst_mult_1_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_107 (
// Equation(s):
// Xd_0__inst_mult_12_340  = SUM(( !Xd_0__inst_mult_12_456  $ (!Xd_0__inst_mult_12_460  $ (Xd_0__inst_mult_12_63_sumout )) ) + ( Xd_0__inst_mult_12_334  ) + ( Xd_0__inst_mult_12_333  ))
// Xd_0__inst_mult_12_341  = CARRY(( !Xd_0__inst_mult_12_456  $ (!Xd_0__inst_mult_12_460  $ (Xd_0__inst_mult_12_63_sumout )) ) + ( Xd_0__inst_mult_12_334  ) + ( Xd_0__inst_mult_12_333  ))
// Xd_0__inst_mult_12_342  = SHARE((!Xd_0__inst_mult_12_456  & (Xd_0__inst_mult_12_460  & Xd_0__inst_mult_12_63_sumout )) # (Xd_0__inst_mult_12_456  & ((Xd_0__inst_mult_12_63_sumout ) # (Xd_0__inst_mult_12_460 ))))

	.dataa(!Xd_0__inst_mult_12_456 ),
	.datab(!Xd_0__inst_mult_12_460 ),
	.datac(!Xd_0__inst_mult_12_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_333 ),
	.sharein(Xd_0__inst_mult_12_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_340 ),
	.cout(Xd_0__inst_mult_12_341 ),
	.shareout(Xd_0__inst_mult_12_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_108 (
// Equation(s):
// Xd_0__inst_mult_12_344  = SUM(( !Xd_0__inst_mult_12_464  $ (((!din_a[145]) # (!din_b[151]))) ) + ( Xd_0__inst_mult_12_470  ) + ( Xd_0__inst_mult_12_469  ))
// Xd_0__inst_mult_12_345  = CARRY(( !Xd_0__inst_mult_12_464  $ (((!din_a[145]) # (!din_b[151]))) ) + ( Xd_0__inst_mult_12_470  ) + ( Xd_0__inst_mult_12_469  ))
// Xd_0__inst_mult_12_346  = SHARE((din_a[145] & (din_b[151] & Xd_0__inst_mult_12_464 )))

	.dataa(!din_a[145]),
	.datab(!din_b[151]),
	.datac(!Xd_0__inst_mult_12_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_469 ),
	.sharein(Xd_0__inst_mult_12_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_344 ),
	.cout(Xd_0__inst_mult_12_345 ),
	.shareout(Xd_0__inst_mult_12_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_105 (
// Equation(s):
// Xd_0__inst_mult_13_320  = SUM(( !Xd_0__inst_mult_13_432  $ (!Xd_0__inst_mult_13_436  $ (Xd_0__inst_mult_13_35_sumout )) ) + ( Xd_0__inst_mult_13_314  ) + ( Xd_0__inst_mult_13_313  ))
// Xd_0__inst_mult_13_321  = CARRY(( !Xd_0__inst_mult_13_432  $ (!Xd_0__inst_mult_13_436  $ (Xd_0__inst_mult_13_35_sumout )) ) + ( Xd_0__inst_mult_13_314  ) + ( Xd_0__inst_mult_13_313  ))
// Xd_0__inst_mult_13_322  = SHARE((!Xd_0__inst_mult_13_432  & (Xd_0__inst_mult_13_436  & Xd_0__inst_mult_13_35_sumout )) # (Xd_0__inst_mult_13_432  & ((Xd_0__inst_mult_13_35_sumout ) # (Xd_0__inst_mult_13_436 ))))

	.dataa(!Xd_0__inst_mult_13_432 ),
	.datab(!Xd_0__inst_mult_13_436 ),
	.datac(!Xd_0__inst_mult_13_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_313 ),
	.sharein(Xd_0__inst_mult_13_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_320 ),
	.cout(Xd_0__inst_mult_13_321 ),
	.shareout(Xd_0__inst_mult_13_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_106 (
// Equation(s):
// Xd_0__inst_mult_13_324  = SUM(( !Xd_0__inst_mult_13_440  $ (((!din_a[157]) # (!din_b[163]))) ) + ( Xd_0__inst_mult_13_446  ) + ( Xd_0__inst_mult_13_445  ))
// Xd_0__inst_mult_13_325  = CARRY(( !Xd_0__inst_mult_13_440  $ (((!din_a[157]) # (!din_b[163]))) ) + ( Xd_0__inst_mult_13_446  ) + ( Xd_0__inst_mult_13_445  ))
// Xd_0__inst_mult_13_326  = SHARE((din_a[157] & (din_b[163] & Xd_0__inst_mult_13_440 )))

	.dataa(!din_a[157]),
	.datab(!din_b[163]),
	.datac(!Xd_0__inst_mult_13_440 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_445 ),
	.sharein(Xd_0__inst_mult_13_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_324 ),
	.cout(Xd_0__inst_mult_13_325 ),
	.shareout(Xd_0__inst_mult_13_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_111 (
// Equation(s):
// Xd_0__inst_mult_14_344  = SUM(( !Xd_0__inst_mult_14_448  $ (!Xd_0__inst_mult_14_452  $ (Xd_0__inst_mult_14_39_sumout )) ) + ( Xd_0__inst_mult_14_338  ) + ( Xd_0__inst_mult_14_337  ))
// Xd_0__inst_mult_14_345  = CARRY(( !Xd_0__inst_mult_14_448  $ (!Xd_0__inst_mult_14_452  $ (Xd_0__inst_mult_14_39_sumout )) ) + ( Xd_0__inst_mult_14_338  ) + ( Xd_0__inst_mult_14_337  ))
// Xd_0__inst_mult_14_346  = SHARE((!Xd_0__inst_mult_14_448  & (Xd_0__inst_mult_14_452  & Xd_0__inst_mult_14_39_sumout )) # (Xd_0__inst_mult_14_448  & ((Xd_0__inst_mult_14_39_sumout ) # (Xd_0__inst_mult_14_452 ))))

	.dataa(!Xd_0__inst_mult_14_448 ),
	.datab(!Xd_0__inst_mult_14_452 ),
	.datac(!Xd_0__inst_mult_14_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_337 ),
	.sharein(Xd_0__inst_mult_14_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_344 ),
	.cout(Xd_0__inst_mult_14_345 ),
	.shareout(Xd_0__inst_mult_14_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_112 (
// Equation(s):
// Xd_0__inst_mult_14_348  = SUM(( !Xd_0__inst_mult_14_456  $ (((!din_a[169]) # (!din_b[175]))) ) + ( Xd_0__inst_mult_14_462  ) + ( Xd_0__inst_mult_14_461  ))
// Xd_0__inst_mult_14_349  = CARRY(( !Xd_0__inst_mult_14_456  $ (((!din_a[169]) # (!din_b[175]))) ) + ( Xd_0__inst_mult_14_462  ) + ( Xd_0__inst_mult_14_461  ))
// Xd_0__inst_mult_14_350  = SHARE((din_a[169] & (din_b[175] & Xd_0__inst_mult_14_456 )))

	.dataa(!din_a[169]),
	.datab(!din_b[175]),
	.datac(!Xd_0__inst_mult_14_456 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_461 ),
	.sharein(Xd_0__inst_mult_14_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_348 ),
	.cout(Xd_0__inst_mult_14_349 ),
	.shareout(Xd_0__inst_mult_14_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_111 (
// Equation(s):
// Xd_0__inst_mult_15_344  = SUM(( !Xd_0__inst_mult_15_460  $ (!Xd_0__inst_mult_15_464  $ (Xd_0__inst_mult_15_43_sumout )) ) + ( Xd_0__inst_mult_15_338  ) + ( Xd_0__inst_mult_15_337  ))
// Xd_0__inst_mult_15_345  = CARRY(( !Xd_0__inst_mult_15_460  $ (!Xd_0__inst_mult_15_464  $ (Xd_0__inst_mult_15_43_sumout )) ) + ( Xd_0__inst_mult_15_338  ) + ( Xd_0__inst_mult_15_337  ))
// Xd_0__inst_mult_15_346  = SHARE((!Xd_0__inst_mult_15_460  & (Xd_0__inst_mult_15_464  & Xd_0__inst_mult_15_43_sumout )) # (Xd_0__inst_mult_15_460  & ((Xd_0__inst_mult_15_43_sumout ) # (Xd_0__inst_mult_15_464 ))))

	.dataa(!Xd_0__inst_mult_15_460 ),
	.datab(!Xd_0__inst_mult_15_464 ),
	.datac(!Xd_0__inst_mult_15_43_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_337 ),
	.sharein(Xd_0__inst_mult_15_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_344 ),
	.cout(Xd_0__inst_mult_15_345 ),
	.shareout(Xd_0__inst_mult_15_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_112 (
// Equation(s):
// Xd_0__inst_mult_15_348  = SUM(( !Xd_0__inst_mult_15_468  $ (((!din_a[181]) # (!din_b[187]))) ) + ( Xd_0__inst_mult_15_474  ) + ( Xd_0__inst_mult_15_473  ))
// Xd_0__inst_mult_15_349  = CARRY(( !Xd_0__inst_mult_15_468  $ (((!din_a[181]) # (!din_b[187]))) ) + ( Xd_0__inst_mult_15_474  ) + ( Xd_0__inst_mult_15_473  ))
// Xd_0__inst_mult_15_350  = SHARE((din_a[181] & (din_b[187] & Xd_0__inst_mult_15_468 )))

	.dataa(!din_a[181]),
	.datab(!din_b[187]),
	.datac(!Xd_0__inst_mult_15_468 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_473 ),
	.sharein(Xd_0__inst_mult_15_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_348 ),
	.cout(Xd_0__inst_mult_15_349 ),
	.shareout(Xd_0__inst_mult_15_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_101 (
// Equation(s):
// Xd_0__inst_mult_10_316  = SUM(( !Xd_0__inst_mult_10_428  $ (!Xd_0__inst_mult_10_432  $ (Xd_0__inst_mult_10_39_sumout )) ) + ( Xd_0__inst_mult_10_310  ) + ( Xd_0__inst_mult_10_309  ))
// Xd_0__inst_mult_10_317  = CARRY(( !Xd_0__inst_mult_10_428  $ (!Xd_0__inst_mult_10_432  $ (Xd_0__inst_mult_10_39_sumout )) ) + ( Xd_0__inst_mult_10_310  ) + ( Xd_0__inst_mult_10_309  ))
// Xd_0__inst_mult_10_318  = SHARE((!Xd_0__inst_mult_10_428  & (Xd_0__inst_mult_10_432  & Xd_0__inst_mult_10_39_sumout )) # (Xd_0__inst_mult_10_428  & ((Xd_0__inst_mult_10_39_sumout ) # (Xd_0__inst_mult_10_432 ))))

	.dataa(!Xd_0__inst_mult_10_428 ),
	.datab(!Xd_0__inst_mult_10_432 ),
	.datac(!Xd_0__inst_mult_10_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_309 ),
	.sharein(Xd_0__inst_mult_10_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_316 ),
	.cout(Xd_0__inst_mult_10_317 ),
	.shareout(Xd_0__inst_mult_10_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_102 (
// Equation(s):
// Xd_0__inst_mult_10_320  = SUM(( !Xd_0__inst_mult_10_436  $ (((!din_a[121]) # (!din_b[127]))) ) + ( Xd_0__inst_mult_10_442  ) + ( Xd_0__inst_mult_10_441  ))
// Xd_0__inst_mult_10_321  = CARRY(( !Xd_0__inst_mult_10_436  $ (((!din_a[121]) # (!din_b[127]))) ) + ( Xd_0__inst_mult_10_442  ) + ( Xd_0__inst_mult_10_441  ))
// Xd_0__inst_mult_10_322  = SHARE((din_a[121] & (din_b[127] & Xd_0__inst_mult_10_436 )))

	.dataa(!din_a[121]),
	.datab(!din_b[127]),
	.datac(!Xd_0__inst_mult_10_436 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_441 ),
	.sharein(Xd_0__inst_mult_10_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_320 ),
	.cout(Xd_0__inst_mult_10_321 ),
	.shareout(Xd_0__inst_mult_10_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_105 (
// Equation(s):
// Xd_0__inst_mult_11_320  = SUM(( !Xd_0__inst_mult_11_432  $ (!Xd_0__inst_mult_11_436  $ (Xd_0__inst_mult_11_59_sumout )) ) + ( Xd_0__inst_mult_11_314  ) + ( Xd_0__inst_mult_11_313  ))
// Xd_0__inst_mult_11_321  = CARRY(( !Xd_0__inst_mult_11_432  $ (!Xd_0__inst_mult_11_436  $ (Xd_0__inst_mult_11_59_sumout )) ) + ( Xd_0__inst_mult_11_314  ) + ( Xd_0__inst_mult_11_313  ))
// Xd_0__inst_mult_11_322  = SHARE((!Xd_0__inst_mult_11_432  & (Xd_0__inst_mult_11_436  & Xd_0__inst_mult_11_59_sumout )) # (Xd_0__inst_mult_11_432  & ((Xd_0__inst_mult_11_59_sumout ) # (Xd_0__inst_mult_11_436 ))))

	.dataa(!Xd_0__inst_mult_11_432 ),
	.datab(!Xd_0__inst_mult_11_436 ),
	.datac(!Xd_0__inst_mult_11_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_313 ),
	.sharein(Xd_0__inst_mult_11_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_320 ),
	.cout(Xd_0__inst_mult_11_321 ),
	.shareout(Xd_0__inst_mult_11_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_106 (
// Equation(s):
// Xd_0__inst_mult_11_324  = SUM(( !Xd_0__inst_mult_11_440  $ (((!din_a[133]) # (!din_b[139]))) ) + ( Xd_0__inst_mult_11_446  ) + ( Xd_0__inst_mult_11_445  ))
// Xd_0__inst_mult_11_325  = CARRY(( !Xd_0__inst_mult_11_440  $ (((!din_a[133]) # (!din_b[139]))) ) + ( Xd_0__inst_mult_11_446  ) + ( Xd_0__inst_mult_11_445  ))
// Xd_0__inst_mult_11_326  = SHARE((din_a[133] & (din_b[139] & Xd_0__inst_mult_11_440 )))

	.dataa(!din_a[133]),
	.datab(!din_b[139]),
	.datac(!Xd_0__inst_mult_11_440 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_445 ),
	.sharein(Xd_0__inst_mult_11_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_324 ),
	.cout(Xd_0__inst_mult_11_325 ),
	.shareout(Xd_0__inst_mult_11_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_105 (
// Equation(s):
// Xd_0__inst_mult_8_320  = SUM(( !Xd_0__inst_mult_8_432  $ (!Xd_0__inst_mult_8_436  $ (Xd_0__inst_mult_8_39_sumout )) ) + ( Xd_0__inst_mult_8_314  ) + ( Xd_0__inst_mult_8_313  ))
// Xd_0__inst_mult_8_321  = CARRY(( !Xd_0__inst_mult_8_432  $ (!Xd_0__inst_mult_8_436  $ (Xd_0__inst_mult_8_39_sumout )) ) + ( Xd_0__inst_mult_8_314  ) + ( Xd_0__inst_mult_8_313  ))
// Xd_0__inst_mult_8_322  = SHARE((!Xd_0__inst_mult_8_432  & (Xd_0__inst_mult_8_436  & Xd_0__inst_mult_8_39_sumout )) # (Xd_0__inst_mult_8_432  & ((Xd_0__inst_mult_8_39_sumout ) # (Xd_0__inst_mult_8_436 ))))

	.dataa(!Xd_0__inst_mult_8_432 ),
	.datab(!Xd_0__inst_mult_8_436 ),
	.datac(!Xd_0__inst_mult_8_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_313 ),
	.sharein(Xd_0__inst_mult_8_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_320 ),
	.cout(Xd_0__inst_mult_8_321 ),
	.shareout(Xd_0__inst_mult_8_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_106 (
// Equation(s):
// Xd_0__inst_mult_8_324  = SUM(( !Xd_0__inst_mult_8_440  $ (((!din_a[97]) # (!din_b[103]))) ) + ( Xd_0__inst_mult_8_446  ) + ( Xd_0__inst_mult_8_445  ))
// Xd_0__inst_mult_8_325  = CARRY(( !Xd_0__inst_mult_8_440  $ (((!din_a[97]) # (!din_b[103]))) ) + ( Xd_0__inst_mult_8_446  ) + ( Xd_0__inst_mult_8_445  ))
// Xd_0__inst_mult_8_326  = SHARE((din_a[97] & (din_b[103] & Xd_0__inst_mult_8_440 )))

	.dataa(!din_a[97]),
	.datab(!din_b[103]),
	.datac(!Xd_0__inst_mult_8_440 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_445 ),
	.sharein(Xd_0__inst_mult_8_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_324 ),
	.cout(Xd_0__inst_mult_8_325 ),
	.shareout(Xd_0__inst_mult_8_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_101 (
// Equation(s):
// Xd_0__inst_mult_9_316  = SUM(( !Xd_0__inst_mult_9_428  $ (!Xd_0__inst_mult_9_432  $ (Xd_0__inst_mult_9_63_sumout )) ) + ( Xd_0__inst_mult_9_310  ) + ( Xd_0__inst_mult_9_309  ))
// Xd_0__inst_mult_9_317  = CARRY(( !Xd_0__inst_mult_9_428  $ (!Xd_0__inst_mult_9_432  $ (Xd_0__inst_mult_9_63_sumout )) ) + ( Xd_0__inst_mult_9_310  ) + ( Xd_0__inst_mult_9_309  ))
// Xd_0__inst_mult_9_318  = SHARE((!Xd_0__inst_mult_9_428  & (Xd_0__inst_mult_9_432  & Xd_0__inst_mult_9_63_sumout )) # (Xd_0__inst_mult_9_428  & ((Xd_0__inst_mult_9_63_sumout ) # (Xd_0__inst_mult_9_432 ))))

	.dataa(!Xd_0__inst_mult_9_428 ),
	.datab(!Xd_0__inst_mult_9_432 ),
	.datac(!Xd_0__inst_mult_9_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_309 ),
	.sharein(Xd_0__inst_mult_9_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_316 ),
	.cout(Xd_0__inst_mult_9_317 ),
	.shareout(Xd_0__inst_mult_9_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_102 (
// Equation(s):
// Xd_0__inst_mult_9_320  = SUM(( !Xd_0__inst_mult_9_436  $ (((!din_a[109]) # (!din_b[115]))) ) + ( Xd_0__inst_mult_9_442  ) + ( Xd_0__inst_mult_9_441  ))
// Xd_0__inst_mult_9_321  = CARRY(( !Xd_0__inst_mult_9_436  $ (((!din_a[109]) # (!din_b[115]))) ) + ( Xd_0__inst_mult_9_442  ) + ( Xd_0__inst_mult_9_441  ))
// Xd_0__inst_mult_9_322  = SHARE((din_a[109] & (din_b[115] & Xd_0__inst_mult_9_436 )))

	.dataa(!din_a[109]),
	.datab(!din_b[115]),
	.datac(!Xd_0__inst_mult_9_436 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_441 ),
	.sharein(Xd_0__inst_mult_9_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_320 ),
	.cout(Xd_0__inst_mult_9_321 ),
	.shareout(Xd_0__inst_mult_9_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_101 (
// Equation(s):
// Xd_0__inst_mult_6_316  = SUM(( !Xd_0__inst_mult_6_428  $ (!Xd_0__inst_mult_6_432  $ (Xd_0__inst_mult_4_420 )) ) + ( Xd_0__inst_mult_6_310  ) + ( Xd_0__inst_mult_6_309  ))
// Xd_0__inst_mult_6_317  = CARRY(( !Xd_0__inst_mult_6_428  $ (!Xd_0__inst_mult_6_432  $ (Xd_0__inst_mult_4_420 )) ) + ( Xd_0__inst_mult_6_310  ) + ( Xd_0__inst_mult_6_309  ))
// Xd_0__inst_mult_6_318  = SHARE((!Xd_0__inst_mult_6_428  & (Xd_0__inst_mult_6_432  & Xd_0__inst_mult_4_420 )) # (Xd_0__inst_mult_6_428  & ((Xd_0__inst_mult_4_420 ) # (Xd_0__inst_mult_6_432 ))))

	.dataa(!Xd_0__inst_mult_6_428 ),
	.datab(!Xd_0__inst_mult_6_432 ),
	.datac(!Xd_0__inst_mult_4_420 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_309 ),
	.sharein(Xd_0__inst_mult_6_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_316 ),
	.cout(Xd_0__inst_mult_6_317 ),
	.shareout(Xd_0__inst_mult_6_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_102 (
// Equation(s):
// Xd_0__inst_mult_6_320  = SUM(( !Xd_0__inst_mult_6_436  $ (((!din_a[73]) # (!din_b[79]))) ) + ( Xd_0__inst_mult_6_442  ) + ( Xd_0__inst_mult_6_441  ))
// Xd_0__inst_mult_6_321  = CARRY(( !Xd_0__inst_mult_6_436  $ (((!din_a[73]) # (!din_b[79]))) ) + ( Xd_0__inst_mult_6_442  ) + ( Xd_0__inst_mult_6_441  ))
// Xd_0__inst_mult_6_322  = SHARE((din_a[73] & (din_b[79] & Xd_0__inst_mult_6_436 )))

	.dataa(!din_a[73]),
	.datab(!din_b[79]),
	.datac(!Xd_0__inst_mult_6_436 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_441 ),
	.sharein(Xd_0__inst_mult_6_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_320 ),
	.cout(Xd_0__inst_mult_6_321 ),
	.shareout(Xd_0__inst_mult_6_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_95 (
// Equation(s):
// Xd_0__inst_mult_7_292  = SUM(( !Xd_0__inst_mult_7_412  $ (!Xd_0__inst_mult_7_416  $ (Xd_0__inst_mult_7_59_sumout )) ) + ( Xd_0__inst_mult_7_286  ) + ( Xd_0__inst_mult_7_285  ))
// Xd_0__inst_mult_7_293  = CARRY(( !Xd_0__inst_mult_7_412  $ (!Xd_0__inst_mult_7_416  $ (Xd_0__inst_mult_7_59_sumout )) ) + ( Xd_0__inst_mult_7_286  ) + ( Xd_0__inst_mult_7_285  ))
// Xd_0__inst_mult_7_294  = SHARE((!Xd_0__inst_mult_7_412  & (Xd_0__inst_mult_7_416  & Xd_0__inst_mult_7_59_sumout )) # (Xd_0__inst_mult_7_412  & ((Xd_0__inst_mult_7_59_sumout ) # (Xd_0__inst_mult_7_416 ))))

	.dataa(!Xd_0__inst_mult_7_412 ),
	.datab(!Xd_0__inst_mult_7_416 ),
	.datac(!Xd_0__inst_mult_7_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_285 ),
	.sharein(Xd_0__inst_mult_7_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_292 ),
	.cout(Xd_0__inst_mult_7_293 ),
	.shareout(Xd_0__inst_mult_7_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_96 (
// Equation(s):
// Xd_0__inst_mult_7_296  = SUM(( !Xd_0__inst_mult_7_420  $ (((!din_a[85]) # (!din_b[91]))) ) + ( Xd_0__inst_mult_7_426  ) + ( Xd_0__inst_mult_7_425  ))
// Xd_0__inst_mult_7_297  = CARRY(( !Xd_0__inst_mult_7_420  $ (((!din_a[85]) # (!din_b[91]))) ) + ( Xd_0__inst_mult_7_426  ) + ( Xd_0__inst_mult_7_425  ))
// Xd_0__inst_mult_7_298  = SHARE((din_a[85] & (din_b[91] & Xd_0__inst_mult_7_420 )))

	.dataa(!din_a[85]),
	.datab(!din_b[91]),
	.datac(!Xd_0__inst_mult_7_420 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_425 ),
	.sharein(Xd_0__inst_mult_7_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_296 ),
	.cout(Xd_0__inst_mult_7_297 ),
	.shareout(Xd_0__inst_mult_7_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_107 (
// Equation(s):
// Xd_0__inst_mult_4_328  = SUM(( !Xd_0__inst_mult_4_452  $ (!Xd_0__inst_mult_4_456  $ (Xd_0__inst_mult_4_63_sumout )) ) + ( Xd_0__inst_mult_4_322  ) + ( Xd_0__inst_mult_4_321  ))
// Xd_0__inst_mult_4_329  = CARRY(( !Xd_0__inst_mult_4_452  $ (!Xd_0__inst_mult_4_456  $ (Xd_0__inst_mult_4_63_sumout )) ) + ( Xd_0__inst_mult_4_322  ) + ( Xd_0__inst_mult_4_321  ))
// Xd_0__inst_mult_4_330  = SHARE((!Xd_0__inst_mult_4_452  & (Xd_0__inst_mult_4_456  & Xd_0__inst_mult_4_63_sumout )) # (Xd_0__inst_mult_4_452  & ((Xd_0__inst_mult_4_63_sumout ) # (Xd_0__inst_mult_4_456 ))))

	.dataa(!Xd_0__inst_mult_4_452 ),
	.datab(!Xd_0__inst_mult_4_456 ),
	.datac(!Xd_0__inst_mult_4_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_321 ),
	.sharein(Xd_0__inst_mult_4_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_328 ),
	.cout(Xd_0__inst_mult_4_329 ),
	.shareout(Xd_0__inst_mult_4_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_108 (
// Equation(s):
// Xd_0__inst_mult_4_332  = SUM(( !Xd_0__inst_mult_4_460  $ (((!din_a[49]) # (!din_b[55]))) ) + ( Xd_0__inst_mult_4_466  ) + ( Xd_0__inst_mult_4_465  ))
// Xd_0__inst_mult_4_333  = CARRY(( !Xd_0__inst_mult_4_460  $ (((!din_a[49]) # (!din_b[55]))) ) + ( Xd_0__inst_mult_4_466  ) + ( Xd_0__inst_mult_4_465  ))
// Xd_0__inst_mult_4_334  = SHARE((din_a[49] & (din_b[55] & Xd_0__inst_mult_4_460 )))

	.dataa(!din_a[49]),
	.datab(!din_b[55]),
	.datac(!Xd_0__inst_mult_4_460 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_465 ),
	.sharein(Xd_0__inst_mult_4_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_332 ),
	.cout(Xd_0__inst_mult_4_333 ),
	.shareout(Xd_0__inst_mult_4_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_95 (
// Equation(s):
// Xd_0__inst_mult_5_292  = SUM(( !Xd_0__inst_mult_5_412  $ (!Xd_0__inst_mult_5_416  $ (Xd_0__inst_mult_5_63_sumout )) ) + ( Xd_0__inst_mult_5_286  ) + ( Xd_0__inst_mult_5_285  ))
// Xd_0__inst_mult_5_293  = CARRY(( !Xd_0__inst_mult_5_412  $ (!Xd_0__inst_mult_5_416  $ (Xd_0__inst_mult_5_63_sumout )) ) + ( Xd_0__inst_mult_5_286  ) + ( Xd_0__inst_mult_5_285  ))
// Xd_0__inst_mult_5_294  = SHARE((!Xd_0__inst_mult_5_412  & (Xd_0__inst_mult_5_416  & Xd_0__inst_mult_5_63_sumout )) # (Xd_0__inst_mult_5_412  & ((Xd_0__inst_mult_5_63_sumout ) # (Xd_0__inst_mult_5_416 ))))

	.dataa(!Xd_0__inst_mult_5_412 ),
	.datab(!Xd_0__inst_mult_5_416 ),
	.datac(!Xd_0__inst_mult_5_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_285 ),
	.sharein(Xd_0__inst_mult_5_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_292 ),
	.cout(Xd_0__inst_mult_5_293 ),
	.shareout(Xd_0__inst_mult_5_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_96 (
// Equation(s):
// Xd_0__inst_mult_5_296  = SUM(( !Xd_0__inst_mult_5_420  $ (((!din_a[61]) # (!din_b[67]))) ) + ( Xd_0__inst_mult_5_426  ) + ( Xd_0__inst_mult_5_425  ))
// Xd_0__inst_mult_5_297  = CARRY(( !Xd_0__inst_mult_5_420  $ (((!din_a[61]) # (!din_b[67]))) ) + ( Xd_0__inst_mult_5_426  ) + ( Xd_0__inst_mult_5_425  ))
// Xd_0__inst_mult_5_298  = SHARE((din_a[61] & (din_b[67] & Xd_0__inst_mult_5_420 )))

	.dataa(!din_a[61]),
	.datab(!din_b[67]),
	.datac(!Xd_0__inst_mult_5_420 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_425 ),
	.sharein(Xd_0__inst_mult_5_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_296 ),
	.cout(Xd_0__inst_mult_5_297 ),
	.shareout(Xd_0__inst_mult_5_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_99 (
// Equation(s):
// Xd_0__inst_mult_2_296  = SUM(( !Xd_0__inst_mult_2_416  $ (!Xd_0__inst_mult_2_420  $ (Xd_0__inst_mult_2_63_sumout )) ) + ( Xd_0__inst_mult_2_290  ) + ( Xd_0__inst_mult_2_289  ))
// Xd_0__inst_mult_2_297  = CARRY(( !Xd_0__inst_mult_2_416  $ (!Xd_0__inst_mult_2_420  $ (Xd_0__inst_mult_2_63_sumout )) ) + ( Xd_0__inst_mult_2_290  ) + ( Xd_0__inst_mult_2_289  ))
// Xd_0__inst_mult_2_298  = SHARE((!Xd_0__inst_mult_2_416  & (Xd_0__inst_mult_2_420  & Xd_0__inst_mult_2_63_sumout )) # (Xd_0__inst_mult_2_416  & ((Xd_0__inst_mult_2_63_sumout ) # (Xd_0__inst_mult_2_420 ))))

	.dataa(!Xd_0__inst_mult_2_416 ),
	.datab(!Xd_0__inst_mult_2_420 ),
	.datac(!Xd_0__inst_mult_2_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_289 ),
	.sharein(Xd_0__inst_mult_2_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_296 ),
	.cout(Xd_0__inst_mult_2_297 ),
	.shareout(Xd_0__inst_mult_2_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_100 (
// Equation(s):
// Xd_0__inst_mult_2_300  = SUM(( !Xd_0__inst_mult_2_424  $ (((!din_a[25]) # (!din_b[31]))) ) + ( Xd_0__inst_mult_2_430  ) + ( Xd_0__inst_mult_2_429  ))
// Xd_0__inst_mult_2_301  = CARRY(( !Xd_0__inst_mult_2_424  $ (((!din_a[25]) # (!din_b[31]))) ) + ( Xd_0__inst_mult_2_430  ) + ( Xd_0__inst_mult_2_429  ))
// Xd_0__inst_mult_2_302  = SHARE((din_a[25] & (din_b[31] & Xd_0__inst_mult_2_424 )))

	.dataa(!din_a[25]),
	.datab(!din_b[31]),
	.datac(!Xd_0__inst_mult_2_424 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_429 ),
	.sharein(Xd_0__inst_mult_2_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_300 ),
	.cout(Xd_0__inst_mult_2_301 ),
	.shareout(Xd_0__inst_mult_2_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_95 (
// Equation(s):
// Xd_0__inst_mult_3_292  = SUM(( !Xd_0__inst_mult_3_412  $ (!Xd_0__inst_mult_3_416  $ (Xd_0__inst_mult_5_380 )) ) + ( Xd_0__inst_mult_3_286  ) + ( Xd_0__inst_mult_3_285  ))
// Xd_0__inst_mult_3_293  = CARRY(( !Xd_0__inst_mult_3_412  $ (!Xd_0__inst_mult_3_416  $ (Xd_0__inst_mult_5_380 )) ) + ( Xd_0__inst_mult_3_286  ) + ( Xd_0__inst_mult_3_285  ))
// Xd_0__inst_mult_3_294  = SHARE((!Xd_0__inst_mult_3_412  & (Xd_0__inst_mult_3_416  & Xd_0__inst_mult_5_380 )) # (Xd_0__inst_mult_3_412  & ((Xd_0__inst_mult_5_380 ) # (Xd_0__inst_mult_3_416 ))))

	.dataa(!Xd_0__inst_mult_3_412 ),
	.datab(!Xd_0__inst_mult_3_416 ),
	.datac(!Xd_0__inst_mult_5_380 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_285 ),
	.sharein(Xd_0__inst_mult_3_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_292 ),
	.cout(Xd_0__inst_mult_3_293 ),
	.shareout(Xd_0__inst_mult_3_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_96 (
// Equation(s):
// Xd_0__inst_mult_3_296  = SUM(( !Xd_0__inst_mult_3_420  $ (((!din_a[37]) # (!din_b[43]))) ) + ( Xd_0__inst_mult_3_426  ) + ( Xd_0__inst_mult_3_425  ))
// Xd_0__inst_mult_3_297  = CARRY(( !Xd_0__inst_mult_3_420  $ (((!din_a[37]) # (!din_b[43]))) ) + ( Xd_0__inst_mult_3_426  ) + ( Xd_0__inst_mult_3_425  ))
// Xd_0__inst_mult_3_298  = SHARE((din_a[37] & (din_b[43] & Xd_0__inst_mult_3_420 )))

	.dataa(!din_a[37]),
	.datab(!din_b[43]),
	.datac(!Xd_0__inst_mult_3_420 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_425 ),
	.sharein(Xd_0__inst_mult_3_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_296 ),
	.cout(Xd_0__inst_mult_3_297 ),
	.shareout(Xd_0__inst_mult_3_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_99 (
// Equation(s):
// Xd_0__inst_mult_0_296  = SUM(( !Xd_0__inst_mult_0_416  $ (!Xd_0__inst_mult_0_420  $ (Xd_0__inst_mult_0_63_sumout )) ) + ( Xd_0__inst_mult_0_290  ) + ( Xd_0__inst_mult_0_289  ))
// Xd_0__inst_mult_0_297  = CARRY(( !Xd_0__inst_mult_0_416  $ (!Xd_0__inst_mult_0_420  $ (Xd_0__inst_mult_0_63_sumout )) ) + ( Xd_0__inst_mult_0_290  ) + ( Xd_0__inst_mult_0_289  ))
// Xd_0__inst_mult_0_298  = SHARE((!Xd_0__inst_mult_0_416  & (Xd_0__inst_mult_0_420  & Xd_0__inst_mult_0_63_sumout )) # (Xd_0__inst_mult_0_416  & ((Xd_0__inst_mult_0_63_sumout ) # (Xd_0__inst_mult_0_420 ))))

	.dataa(!Xd_0__inst_mult_0_416 ),
	.datab(!Xd_0__inst_mult_0_420 ),
	.datac(!Xd_0__inst_mult_0_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_289 ),
	.sharein(Xd_0__inst_mult_0_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_296 ),
	.cout(Xd_0__inst_mult_0_297 ),
	.shareout(Xd_0__inst_mult_0_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_100 (
// Equation(s):
// Xd_0__inst_mult_0_300  = SUM(( !Xd_0__inst_mult_0_424  $ (((!din_a[1]) # (!din_b[7]))) ) + ( Xd_0__inst_mult_0_430  ) + ( Xd_0__inst_mult_0_429  ))
// Xd_0__inst_mult_0_301  = CARRY(( !Xd_0__inst_mult_0_424  $ (((!din_a[1]) # (!din_b[7]))) ) + ( Xd_0__inst_mult_0_430  ) + ( Xd_0__inst_mult_0_429  ))
// Xd_0__inst_mult_0_302  = SHARE((din_a[1] & (din_b[7] & Xd_0__inst_mult_0_424 )))

	.dataa(!din_a[1]),
	.datab(!din_b[7]),
	.datac(!Xd_0__inst_mult_0_424 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_429 ),
	.sharein(Xd_0__inst_mult_0_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_300 ),
	.cout(Xd_0__inst_mult_0_301 ),
	.shareout(Xd_0__inst_mult_0_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_99 (
// Equation(s):
// Xd_0__inst_mult_1_296  = SUM(( !Xd_0__inst_mult_1_416  $ (!Xd_0__inst_mult_1_420  $ (Xd_0__inst_mult_1_67_sumout )) ) + ( Xd_0__inst_mult_1_290  ) + ( Xd_0__inst_mult_1_289  ))
// Xd_0__inst_mult_1_297  = CARRY(( !Xd_0__inst_mult_1_416  $ (!Xd_0__inst_mult_1_420  $ (Xd_0__inst_mult_1_67_sumout )) ) + ( Xd_0__inst_mult_1_290  ) + ( Xd_0__inst_mult_1_289  ))
// Xd_0__inst_mult_1_298  = SHARE((!Xd_0__inst_mult_1_416  & (Xd_0__inst_mult_1_420  & Xd_0__inst_mult_1_67_sumout )) # (Xd_0__inst_mult_1_416  & ((Xd_0__inst_mult_1_67_sumout ) # (Xd_0__inst_mult_1_420 ))))

	.dataa(!Xd_0__inst_mult_1_416 ),
	.datab(!Xd_0__inst_mult_1_420 ),
	.datac(!Xd_0__inst_mult_1_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_289 ),
	.sharein(Xd_0__inst_mult_1_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_296 ),
	.cout(Xd_0__inst_mult_1_297 ),
	.shareout(Xd_0__inst_mult_1_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_100 (
// Equation(s):
// Xd_0__inst_mult_1_300  = SUM(( !Xd_0__inst_mult_1_424  $ (((!din_a[13]) # (!din_b[19]))) ) + ( Xd_0__inst_mult_1_430  ) + ( Xd_0__inst_mult_1_429  ))
// Xd_0__inst_mult_1_301  = CARRY(( !Xd_0__inst_mult_1_424  $ (((!din_a[13]) # (!din_b[19]))) ) + ( Xd_0__inst_mult_1_430  ) + ( Xd_0__inst_mult_1_429  ))
// Xd_0__inst_mult_1_302  = SHARE((din_a[13] & (din_b[19] & Xd_0__inst_mult_1_424 )))

	.dataa(!din_a[13]),
	.datab(!din_b[19]),
	.datac(!Xd_0__inst_mult_1_424 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_429 ),
	.sharein(Xd_0__inst_mult_1_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_300 ),
	.cout(Xd_0__inst_mult_1_301 ),
	.shareout(Xd_0__inst_mult_1_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_109 (
// Equation(s):
// Xd_0__inst_mult_12_348  = SUM(( !Xd_0__inst_mult_12_472  $ (!Xd_0__inst_mult_12_476  $ (Xd_0__inst_mult_2_384 )) ) + ( Xd_0__inst_mult_12_342  ) + ( Xd_0__inst_mult_12_341  ))
// Xd_0__inst_mult_12_349  = CARRY(( !Xd_0__inst_mult_12_472  $ (!Xd_0__inst_mult_12_476  $ (Xd_0__inst_mult_2_384 )) ) + ( Xd_0__inst_mult_12_342  ) + ( Xd_0__inst_mult_12_341  ))
// Xd_0__inst_mult_12_350  = SHARE((!Xd_0__inst_mult_12_472  & (Xd_0__inst_mult_12_476  & Xd_0__inst_mult_2_384 )) # (Xd_0__inst_mult_12_472  & ((Xd_0__inst_mult_2_384 ) # (Xd_0__inst_mult_12_476 ))))

	.dataa(!Xd_0__inst_mult_12_472 ),
	.datab(!Xd_0__inst_mult_12_476 ),
	.datac(!Xd_0__inst_mult_2_384 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_341 ),
	.sharein(Xd_0__inst_mult_12_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_348 ),
	.cout(Xd_0__inst_mult_12_349 ),
	.shareout(Xd_0__inst_mult_12_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_110 (
// Equation(s):
// Xd_0__inst_mult_12_352  = SUM(( !Xd_0__inst_mult_12_480  $ (!Xd_0__inst_mult_12_484 ) ) + ( Xd_0__inst_mult_12_346  ) + ( Xd_0__inst_mult_12_345  ))
// Xd_0__inst_mult_12_353  = CARRY(( !Xd_0__inst_mult_12_480  $ (!Xd_0__inst_mult_12_484 ) ) + ( Xd_0__inst_mult_12_346  ) + ( Xd_0__inst_mult_12_345  ))
// Xd_0__inst_mult_12_354  = SHARE((Xd_0__inst_mult_12_480  & Xd_0__inst_mult_12_484 ))

	.dataa(!Xd_0__inst_mult_12_480 ),
	.datab(!Xd_0__inst_mult_12_484 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_345 ),
	.sharein(Xd_0__inst_mult_12_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_352 ),
	.cout(Xd_0__inst_mult_12_353 ),
	.shareout(Xd_0__inst_mult_12_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_107 (
// Equation(s):
// Xd_0__inst_mult_13_328  = SUM(( !Xd_0__inst_mult_13_448  $ (!Xd_0__inst_mult_13_452  $ (Xd_0__inst_mult_13_67_sumout )) ) + ( Xd_0__inst_mult_13_322  ) + ( Xd_0__inst_mult_13_321  ))
// Xd_0__inst_mult_13_329  = CARRY(( !Xd_0__inst_mult_13_448  $ (!Xd_0__inst_mult_13_452  $ (Xd_0__inst_mult_13_67_sumout )) ) + ( Xd_0__inst_mult_13_322  ) + ( Xd_0__inst_mult_13_321  ))
// Xd_0__inst_mult_13_330  = SHARE((!Xd_0__inst_mult_13_448  & (Xd_0__inst_mult_13_452  & Xd_0__inst_mult_13_67_sumout )) # (Xd_0__inst_mult_13_448  & ((Xd_0__inst_mult_13_67_sumout ) # (Xd_0__inst_mult_13_452 ))))

	.dataa(!Xd_0__inst_mult_13_448 ),
	.datab(!Xd_0__inst_mult_13_452 ),
	.datac(!Xd_0__inst_mult_13_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_321 ),
	.sharein(Xd_0__inst_mult_13_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_328 ),
	.cout(Xd_0__inst_mult_13_329 ),
	.shareout(Xd_0__inst_mult_13_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_108 (
// Equation(s):
// Xd_0__inst_mult_13_332  = SUM(( !Xd_0__inst_mult_13_456  $ (!Xd_0__inst_mult_13_460 ) ) + ( Xd_0__inst_mult_13_326  ) + ( Xd_0__inst_mult_13_325  ))
// Xd_0__inst_mult_13_333  = CARRY(( !Xd_0__inst_mult_13_456  $ (!Xd_0__inst_mult_13_460 ) ) + ( Xd_0__inst_mult_13_326  ) + ( Xd_0__inst_mult_13_325  ))
// Xd_0__inst_mult_13_334  = SHARE((Xd_0__inst_mult_13_456  & Xd_0__inst_mult_13_460 ))

	.dataa(!Xd_0__inst_mult_13_456 ),
	.datab(!Xd_0__inst_mult_13_460 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_325 ),
	.sharein(Xd_0__inst_mult_13_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_332 ),
	.cout(Xd_0__inst_mult_13_333 ),
	.shareout(Xd_0__inst_mult_13_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_113 (
// Equation(s):
// Xd_0__inst_mult_14_352  = SUM(( !Xd_0__inst_mult_14_464  $ (!Xd_0__inst_mult_14_468  $ (Xd_0__inst_mult_14_67_sumout )) ) + ( Xd_0__inst_mult_14_346  ) + ( Xd_0__inst_mult_14_345  ))
// Xd_0__inst_mult_14_353  = CARRY(( !Xd_0__inst_mult_14_464  $ (!Xd_0__inst_mult_14_468  $ (Xd_0__inst_mult_14_67_sumout )) ) + ( Xd_0__inst_mult_14_346  ) + ( Xd_0__inst_mult_14_345  ))
// Xd_0__inst_mult_14_354  = SHARE((!Xd_0__inst_mult_14_464  & (Xd_0__inst_mult_14_468  & Xd_0__inst_mult_14_67_sumout )) # (Xd_0__inst_mult_14_464  & ((Xd_0__inst_mult_14_67_sumout ) # (Xd_0__inst_mult_14_468 ))))

	.dataa(!Xd_0__inst_mult_14_464 ),
	.datab(!Xd_0__inst_mult_14_468 ),
	.datac(!Xd_0__inst_mult_14_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_345 ),
	.sharein(Xd_0__inst_mult_14_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_352 ),
	.cout(Xd_0__inst_mult_14_353 ),
	.shareout(Xd_0__inst_mult_14_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_114 (
// Equation(s):
// Xd_0__inst_mult_14_356  = SUM(( !Xd_0__inst_mult_14_472  $ (!Xd_0__inst_mult_14_476 ) ) + ( Xd_0__inst_mult_14_350  ) + ( Xd_0__inst_mult_14_349  ))
// Xd_0__inst_mult_14_357  = CARRY(( !Xd_0__inst_mult_14_472  $ (!Xd_0__inst_mult_14_476 ) ) + ( Xd_0__inst_mult_14_350  ) + ( Xd_0__inst_mult_14_349  ))
// Xd_0__inst_mult_14_358  = SHARE((Xd_0__inst_mult_14_472  & Xd_0__inst_mult_14_476 ))

	.dataa(!Xd_0__inst_mult_14_472 ),
	.datab(!Xd_0__inst_mult_14_476 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_349 ),
	.sharein(Xd_0__inst_mult_14_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_356 ),
	.cout(Xd_0__inst_mult_14_357 ),
	.shareout(Xd_0__inst_mult_14_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_113 (
// Equation(s):
// Xd_0__inst_mult_15_352  = SUM(( !Xd_0__inst_mult_15_476  $ (!Xd_0__inst_mult_15_480  $ (Xd_0__inst_mult_15_67_sumout )) ) + ( Xd_0__inst_mult_15_346  ) + ( Xd_0__inst_mult_15_345  ))
// Xd_0__inst_mult_15_353  = CARRY(( !Xd_0__inst_mult_15_476  $ (!Xd_0__inst_mult_15_480  $ (Xd_0__inst_mult_15_67_sumout )) ) + ( Xd_0__inst_mult_15_346  ) + ( Xd_0__inst_mult_15_345  ))
// Xd_0__inst_mult_15_354  = SHARE((!Xd_0__inst_mult_15_476  & (Xd_0__inst_mult_15_480  & Xd_0__inst_mult_15_67_sumout )) # (Xd_0__inst_mult_15_476  & ((Xd_0__inst_mult_15_67_sumout ) # (Xd_0__inst_mult_15_480 ))))

	.dataa(!Xd_0__inst_mult_15_476 ),
	.datab(!Xd_0__inst_mult_15_480 ),
	.datac(!Xd_0__inst_mult_15_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_345 ),
	.sharein(Xd_0__inst_mult_15_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_352 ),
	.cout(Xd_0__inst_mult_15_353 ),
	.shareout(Xd_0__inst_mult_15_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_114 (
// Equation(s):
// Xd_0__inst_mult_15_356  = SUM(( !Xd_0__inst_mult_15_484  $ (!Xd_0__inst_mult_15_488 ) ) + ( Xd_0__inst_mult_15_350  ) + ( Xd_0__inst_mult_15_349  ))
// Xd_0__inst_mult_15_357  = CARRY(( !Xd_0__inst_mult_15_484  $ (!Xd_0__inst_mult_15_488 ) ) + ( Xd_0__inst_mult_15_350  ) + ( Xd_0__inst_mult_15_349  ))
// Xd_0__inst_mult_15_358  = SHARE((Xd_0__inst_mult_15_484  & Xd_0__inst_mult_15_488 ))

	.dataa(!Xd_0__inst_mult_15_484 ),
	.datab(!Xd_0__inst_mult_15_488 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_349 ),
	.sharein(Xd_0__inst_mult_15_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_356 ),
	.cout(Xd_0__inst_mult_15_357 ),
	.shareout(Xd_0__inst_mult_15_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_103 (
// Equation(s):
// Xd_0__inst_mult_10_324  = SUM(( !Xd_0__inst_mult_10_444  $ (!Xd_0__inst_mult_10_448  $ (Xd_0__inst_mult_10_63_sumout )) ) + ( Xd_0__inst_mult_10_318  ) + ( Xd_0__inst_mult_10_317  ))
// Xd_0__inst_mult_10_325  = CARRY(( !Xd_0__inst_mult_10_444  $ (!Xd_0__inst_mult_10_448  $ (Xd_0__inst_mult_10_63_sumout )) ) + ( Xd_0__inst_mult_10_318  ) + ( Xd_0__inst_mult_10_317  ))
// Xd_0__inst_mult_10_326  = SHARE((!Xd_0__inst_mult_10_444  & (Xd_0__inst_mult_10_448  & Xd_0__inst_mult_10_63_sumout )) # (Xd_0__inst_mult_10_444  & ((Xd_0__inst_mult_10_63_sumout ) # (Xd_0__inst_mult_10_448 ))))

	.dataa(!Xd_0__inst_mult_10_444 ),
	.datab(!Xd_0__inst_mult_10_448 ),
	.datac(!Xd_0__inst_mult_10_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_317 ),
	.sharein(Xd_0__inst_mult_10_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_324 ),
	.cout(Xd_0__inst_mult_10_325 ),
	.shareout(Xd_0__inst_mult_10_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_104 (
// Equation(s):
// Xd_0__inst_mult_10_328  = SUM(( !Xd_0__inst_mult_10_452  $ (!Xd_0__inst_mult_10_456 ) ) + ( Xd_0__inst_mult_10_322  ) + ( Xd_0__inst_mult_10_321  ))
// Xd_0__inst_mult_10_329  = CARRY(( !Xd_0__inst_mult_10_452  $ (!Xd_0__inst_mult_10_456 ) ) + ( Xd_0__inst_mult_10_322  ) + ( Xd_0__inst_mult_10_321  ))
// Xd_0__inst_mult_10_330  = SHARE((Xd_0__inst_mult_10_452  & Xd_0__inst_mult_10_456 ))

	.dataa(!Xd_0__inst_mult_10_452 ),
	.datab(!Xd_0__inst_mult_10_456 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_321 ),
	.sharein(Xd_0__inst_mult_10_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_328 ),
	.cout(Xd_0__inst_mult_10_329 ),
	.shareout(Xd_0__inst_mult_10_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_107 (
// Equation(s):
// Xd_0__inst_mult_11_328  = SUM(( !Xd_0__inst_mult_11_448  $ (!Xd_0__inst_mult_11_452  $ (Xd_0__inst_mult_11_67_sumout )) ) + ( Xd_0__inst_mult_11_322  ) + ( Xd_0__inst_mult_11_321  ))
// Xd_0__inst_mult_11_329  = CARRY(( !Xd_0__inst_mult_11_448  $ (!Xd_0__inst_mult_11_452  $ (Xd_0__inst_mult_11_67_sumout )) ) + ( Xd_0__inst_mult_11_322  ) + ( Xd_0__inst_mult_11_321  ))
// Xd_0__inst_mult_11_330  = SHARE((!Xd_0__inst_mult_11_448  & (Xd_0__inst_mult_11_452  & Xd_0__inst_mult_11_67_sumout )) # (Xd_0__inst_mult_11_448  & ((Xd_0__inst_mult_11_67_sumout ) # (Xd_0__inst_mult_11_452 ))))

	.dataa(!Xd_0__inst_mult_11_448 ),
	.datab(!Xd_0__inst_mult_11_452 ),
	.datac(!Xd_0__inst_mult_11_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_321 ),
	.sharein(Xd_0__inst_mult_11_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_328 ),
	.cout(Xd_0__inst_mult_11_329 ),
	.shareout(Xd_0__inst_mult_11_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_108 (
// Equation(s):
// Xd_0__inst_mult_11_332  = SUM(( !Xd_0__inst_mult_11_456  $ (!Xd_0__inst_mult_11_460 ) ) + ( Xd_0__inst_mult_11_326  ) + ( Xd_0__inst_mult_11_325  ))
// Xd_0__inst_mult_11_333  = CARRY(( !Xd_0__inst_mult_11_456  $ (!Xd_0__inst_mult_11_460 ) ) + ( Xd_0__inst_mult_11_326  ) + ( Xd_0__inst_mult_11_325  ))
// Xd_0__inst_mult_11_334  = SHARE((Xd_0__inst_mult_11_456  & Xd_0__inst_mult_11_460 ))

	.dataa(!Xd_0__inst_mult_11_456 ),
	.datab(!Xd_0__inst_mult_11_460 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_325 ),
	.sharein(Xd_0__inst_mult_11_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_332 ),
	.cout(Xd_0__inst_mult_11_333 ),
	.shareout(Xd_0__inst_mult_11_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_107 (
// Equation(s):
// Xd_0__inst_mult_8_328  = SUM(( !Xd_0__inst_mult_8_448  $ (!Xd_0__inst_mult_8_452  $ (Xd_0__inst_mult_8_67_sumout )) ) + ( Xd_0__inst_mult_8_322  ) + ( Xd_0__inst_mult_8_321  ))
// Xd_0__inst_mult_8_329  = CARRY(( !Xd_0__inst_mult_8_448  $ (!Xd_0__inst_mult_8_452  $ (Xd_0__inst_mult_8_67_sumout )) ) + ( Xd_0__inst_mult_8_322  ) + ( Xd_0__inst_mult_8_321  ))
// Xd_0__inst_mult_8_330  = SHARE((!Xd_0__inst_mult_8_448  & (Xd_0__inst_mult_8_452  & Xd_0__inst_mult_8_67_sumout )) # (Xd_0__inst_mult_8_448  & ((Xd_0__inst_mult_8_67_sumout ) # (Xd_0__inst_mult_8_452 ))))

	.dataa(!Xd_0__inst_mult_8_448 ),
	.datab(!Xd_0__inst_mult_8_452 ),
	.datac(!Xd_0__inst_mult_8_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_321 ),
	.sharein(Xd_0__inst_mult_8_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_328 ),
	.cout(Xd_0__inst_mult_8_329 ),
	.shareout(Xd_0__inst_mult_8_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_108 (
// Equation(s):
// Xd_0__inst_mult_8_332  = SUM(( !Xd_0__inst_mult_8_456  $ (!Xd_0__inst_mult_8_460 ) ) + ( Xd_0__inst_mult_8_326  ) + ( Xd_0__inst_mult_8_325  ))
// Xd_0__inst_mult_8_333  = CARRY(( !Xd_0__inst_mult_8_456  $ (!Xd_0__inst_mult_8_460 ) ) + ( Xd_0__inst_mult_8_326  ) + ( Xd_0__inst_mult_8_325  ))
// Xd_0__inst_mult_8_334  = SHARE((Xd_0__inst_mult_8_456  & Xd_0__inst_mult_8_460 ))

	.dataa(!Xd_0__inst_mult_8_456 ),
	.datab(!Xd_0__inst_mult_8_460 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_325 ),
	.sharein(Xd_0__inst_mult_8_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_332 ),
	.cout(Xd_0__inst_mult_8_333 ),
	.shareout(Xd_0__inst_mult_8_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_103 (
// Equation(s):
// Xd_0__inst_mult_9_324  = SUM(( !Xd_0__inst_mult_9_444  $ (!Xd_0__inst_mult_9_448  $ (Xd_0__inst_mult_3_380 )) ) + ( Xd_0__inst_mult_9_318  ) + ( Xd_0__inst_mult_9_317  ))
// Xd_0__inst_mult_9_325  = CARRY(( !Xd_0__inst_mult_9_444  $ (!Xd_0__inst_mult_9_448  $ (Xd_0__inst_mult_3_380 )) ) + ( Xd_0__inst_mult_9_318  ) + ( Xd_0__inst_mult_9_317  ))
// Xd_0__inst_mult_9_326  = SHARE((!Xd_0__inst_mult_9_444  & (Xd_0__inst_mult_9_448  & Xd_0__inst_mult_3_380 )) # (Xd_0__inst_mult_9_444  & ((Xd_0__inst_mult_3_380 ) # (Xd_0__inst_mult_9_448 ))))

	.dataa(!Xd_0__inst_mult_9_444 ),
	.datab(!Xd_0__inst_mult_9_448 ),
	.datac(!Xd_0__inst_mult_3_380 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_317 ),
	.sharein(Xd_0__inst_mult_9_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_324 ),
	.cout(Xd_0__inst_mult_9_325 ),
	.shareout(Xd_0__inst_mult_9_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_104 (
// Equation(s):
// Xd_0__inst_mult_9_328  = SUM(( !Xd_0__inst_mult_9_452  $ (!Xd_0__inst_mult_9_456 ) ) + ( Xd_0__inst_mult_9_322  ) + ( Xd_0__inst_mult_9_321  ))
// Xd_0__inst_mult_9_329  = CARRY(( !Xd_0__inst_mult_9_452  $ (!Xd_0__inst_mult_9_456 ) ) + ( Xd_0__inst_mult_9_322  ) + ( Xd_0__inst_mult_9_321  ))
// Xd_0__inst_mult_9_330  = SHARE((Xd_0__inst_mult_9_452  & Xd_0__inst_mult_9_456 ))

	.dataa(!Xd_0__inst_mult_9_452 ),
	.datab(!Xd_0__inst_mult_9_456 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_321 ),
	.sharein(Xd_0__inst_mult_9_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_328 ),
	.cout(Xd_0__inst_mult_9_329 ),
	.shareout(Xd_0__inst_mult_9_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_103 (
// Equation(s):
// Xd_0__inst_mult_6_324  = SUM(( !Xd_0__inst_mult_6_444  $ (!Xd_0__inst_mult_6_448  $ (Xd_0__inst_mult_6_63_sumout )) ) + ( Xd_0__inst_mult_6_318  ) + ( Xd_0__inst_mult_6_317  ))
// Xd_0__inst_mult_6_325  = CARRY(( !Xd_0__inst_mult_6_444  $ (!Xd_0__inst_mult_6_448  $ (Xd_0__inst_mult_6_63_sumout )) ) + ( Xd_0__inst_mult_6_318  ) + ( Xd_0__inst_mult_6_317  ))
// Xd_0__inst_mult_6_326  = SHARE((!Xd_0__inst_mult_6_444  & (Xd_0__inst_mult_6_448  & Xd_0__inst_mult_6_63_sumout )) # (Xd_0__inst_mult_6_444  & ((Xd_0__inst_mult_6_63_sumout ) # (Xd_0__inst_mult_6_448 ))))

	.dataa(!Xd_0__inst_mult_6_444 ),
	.datab(!Xd_0__inst_mult_6_448 ),
	.datac(!Xd_0__inst_mult_6_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_317 ),
	.sharein(Xd_0__inst_mult_6_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_324 ),
	.cout(Xd_0__inst_mult_6_325 ),
	.shareout(Xd_0__inst_mult_6_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_104 (
// Equation(s):
// Xd_0__inst_mult_6_328  = SUM(( !Xd_0__inst_mult_6_452  $ (!Xd_0__inst_mult_6_456 ) ) + ( Xd_0__inst_mult_6_322  ) + ( Xd_0__inst_mult_6_321  ))
// Xd_0__inst_mult_6_329  = CARRY(( !Xd_0__inst_mult_6_452  $ (!Xd_0__inst_mult_6_456 ) ) + ( Xd_0__inst_mult_6_322  ) + ( Xd_0__inst_mult_6_321  ))
// Xd_0__inst_mult_6_330  = SHARE((Xd_0__inst_mult_6_452  & Xd_0__inst_mult_6_456 ))

	.dataa(!Xd_0__inst_mult_6_452 ),
	.datab(!Xd_0__inst_mult_6_456 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_321 ),
	.sharein(Xd_0__inst_mult_6_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_328 ),
	.cout(Xd_0__inst_mult_6_329 ),
	.shareout(Xd_0__inst_mult_6_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_97 (
// Equation(s):
// Xd_0__inst_mult_7_300  = SUM(( !Xd_0__inst_mult_7_428  $ (!Xd_0__inst_mult_7_432  $ (Xd_0__inst_mult_7_63_sumout )) ) + ( Xd_0__inst_mult_7_294  ) + ( Xd_0__inst_mult_7_293  ))
// Xd_0__inst_mult_7_301  = CARRY(( !Xd_0__inst_mult_7_428  $ (!Xd_0__inst_mult_7_432  $ (Xd_0__inst_mult_7_63_sumout )) ) + ( Xd_0__inst_mult_7_294  ) + ( Xd_0__inst_mult_7_293  ))
// Xd_0__inst_mult_7_302  = SHARE((!Xd_0__inst_mult_7_428  & (Xd_0__inst_mult_7_432  & Xd_0__inst_mult_7_63_sumout )) # (Xd_0__inst_mult_7_428  & ((Xd_0__inst_mult_7_63_sumout ) # (Xd_0__inst_mult_7_432 ))))

	.dataa(!Xd_0__inst_mult_7_428 ),
	.datab(!Xd_0__inst_mult_7_432 ),
	.datac(!Xd_0__inst_mult_7_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_293 ),
	.sharein(Xd_0__inst_mult_7_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_300 ),
	.cout(Xd_0__inst_mult_7_301 ),
	.shareout(Xd_0__inst_mult_7_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_98 (
// Equation(s):
// Xd_0__inst_mult_7_304  = SUM(( !Xd_0__inst_mult_7_436  $ (!Xd_0__inst_mult_7_440 ) ) + ( Xd_0__inst_mult_7_298  ) + ( Xd_0__inst_mult_7_297  ))
// Xd_0__inst_mult_7_305  = CARRY(( !Xd_0__inst_mult_7_436  $ (!Xd_0__inst_mult_7_440 ) ) + ( Xd_0__inst_mult_7_298  ) + ( Xd_0__inst_mult_7_297  ))
// Xd_0__inst_mult_7_306  = SHARE((Xd_0__inst_mult_7_436  & Xd_0__inst_mult_7_440 ))

	.dataa(!Xd_0__inst_mult_7_436 ),
	.datab(!Xd_0__inst_mult_7_440 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_297 ),
	.sharein(Xd_0__inst_mult_7_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_304 ),
	.cout(Xd_0__inst_mult_7_305 ),
	.shareout(Xd_0__inst_mult_7_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_109 (
// Equation(s):
// Xd_0__inst_mult_4_336  = SUM(( !Xd_0__inst_mult_4_468  $ (!Xd_0__inst_mult_4_472  $ (Xd_0__inst_mult_4_67_sumout )) ) + ( Xd_0__inst_mult_4_330  ) + ( Xd_0__inst_mult_4_329  ))
// Xd_0__inst_mult_4_337  = CARRY(( !Xd_0__inst_mult_4_468  $ (!Xd_0__inst_mult_4_472  $ (Xd_0__inst_mult_4_67_sumout )) ) + ( Xd_0__inst_mult_4_330  ) + ( Xd_0__inst_mult_4_329  ))
// Xd_0__inst_mult_4_338  = SHARE((!Xd_0__inst_mult_4_468  & (Xd_0__inst_mult_4_472  & Xd_0__inst_mult_4_67_sumout )) # (Xd_0__inst_mult_4_468  & ((Xd_0__inst_mult_4_67_sumout ) # (Xd_0__inst_mult_4_472 ))))

	.dataa(!Xd_0__inst_mult_4_468 ),
	.datab(!Xd_0__inst_mult_4_472 ),
	.datac(!Xd_0__inst_mult_4_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_329 ),
	.sharein(Xd_0__inst_mult_4_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_336 ),
	.cout(Xd_0__inst_mult_4_337 ),
	.shareout(Xd_0__inst_mult_4_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_110 (
// Equation(s):
// Xd_0__inst_mult_4_340  = SUM(( !Xd_0__inst_mult_4_476  $ (!Xd_0__inst_mult_4_480 ) ) + ( Xd_0__inst_mult_4_334  ) + ( Xd_0__inst_mult_4_333  ))
// Xd_0__inst_mult_4_341  = CARRY(( !Xd_0__inst_mult_4_476  $ (!Xd_0__inst_mult_4_480 ) ) + ( Xd_0__inst_mult_4_334  ) + ( Xd_0__inst_mult_4_333  ))
// Xd_0__inst_mult_4_342  = SHARE((Xd_0__inst_mult_4_476  & Xd_0__inst_mult_4_480 ))

	.dataa(!Xd_0__inst_mult_4_476 ),
	.datab(!Xd_0__inst_mult_4_480 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_333 ),
	.sharein(Xd_0__inst_mult_4_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_340 ),
	.cout(Xd_0__inst_mult_4_341 ),
	.shareout(Xd_0__inst_mult_4_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_97 (
// Equation(s):
// Xd_0__inst_mult_5_300  = SUM(( !Xd_0__inst_mult_5_428  $ (!Xd_0__inst_mult_5_432  $ (Xd_0__inst_mult_5_35_sumout )) ) + ( Xd_0__inst_mult_5_294  ) + ( Xd_0__inst_mult_5_293  ))
// Xd_0__inst_mult_5_301  = CARRY(( !Xd_0__inst_mult_5_428  $ (!Xd_0__inst_mult_5_432  $ (Xd_0__inst_mult_5_35_sumout )) ) + ( Xd_0__inst_mult_5_294  ) + ( Xd_0__inst_mult_5_293  ))
// Xd_0__inst_mult_5_302  = SHARE((!Xd_0__inst_mult_5_428  & (Xd_0__inst_mult_5_432  & Xd_0__inst_mult_5_35_sumout )) # (Xd_0__inst_mult_5_428  & ((Xd_0__inst_mult_5_35_sumout ) # (Xd_0__inst_mult_5_432 ))))

	.dataa(!Xd_0__inst_mult_5_428 ),
	.datab(!Xd_0__inst_mult_5_432 ),
	.datac(!Xd_0__inst_mult_5_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_293 ),
	.sharein(Xd_0__inst_mult_5_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_300 ),
	.cout(Xd_0__inst_mult_5_301 ),
	.shareout(Xd_0__inst_mult_5_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_98 (
// Equation(s):
// Xd_0__inst_mult_5_304  = SUM(( !Xd_0__inst_mult_5_436  $ (!Xd_0__inst_mult_5_440 ) ) + ( Xd_0__inst_mult_5_298  ) + ( Xd_0__inst_mult_5_297  ))
// Xd_0__inst_mult_5_305  = CARRY(( !Xd_0__inst_mult_5_436  $ (!Xd_0__inst_mult_5_440 ) ) + ( Xd_0__inst_mult_5_298  ) + ( Xd_0__inst_mult_5_297  ))
// Xd_0__inst_mult_5_306  = SHARE((Xd_0__inst_mult_5_436  & Xd_0__inst_mult_5_440 ))

	.dataa(!Xd_0__inst_mult_5_436 ),
	.datab(!Xd_0__inst_mult_5_440 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_297 ),
	.sharein(Xd_0__inst_mult_5_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_304 ),
	.cout(Xd_0__inst_mult_5_305 ),
	.shareout(Xd_0__inst_mult_5_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_101 (
// Equation(s):
// Xd_0__inst_mult_2_304  = SUM(( !Xd_0__inst_mult_2_432  $ (!Xd_0__inst_mult_2_436  $ (Xd_0__inst_mult_2_35_sumout )) ) + ( Xd_0__inst_mult_2_298  ) + ( Xd_0__inst_mult_2_297  ))
// Xd_0__inst_mult_2_305  = CARRY(( !Xd_0__inst_mult_2_432  $ (!Xd_0__inst_mult_2_436  $ (Xd_0__inst_mult_2_35_sumout )) ) + ( Xd_0__inst_mult_2_298  ) + ( Xd_0__inst_mult_2_297  ))
// Xd_0__inst_mult_2_306  = SHARE((!Xd_0__inst_mult_2_432  & (Xd_0__inst_mult_2_436  & Xd_0__inst_mult_2_35_sumout )) # (Xd_0__inst_mult_2_432  & ((Xd_0__inst_mult_2_35_sumout ) # (Xd_0__inst_mult_2_436 ))))

	.dataa(!Xd_0__inst_mult_2_432 ),
	.datab(!Xd_0__inst_mult_2_436 ),
	.datac(!Xd_0__inst_mult_2_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_297 ),
	.sharein(Xd_0__inst_mult_2_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_304 ),
	.cout(Xd_0__inst_mult_2_305 ),
	.shareout(Xd_0__inst_mult_2_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_102 (
// Equation(s):
// Xd_0__inst_mult_2_308  = SUM(( !Xd_0__inst_mult_2_440  $ (!Xd_0__inst_mult_2_444 ) ) + ( Xd_0__inst_mult_2_302  ) + ( Xd_0__inst_mult_2_301  ))
// Xd_0__inst_mult_2_309  = CARRY(( !Xd_0__inst_mult_2_440  $ (!Xd_0__inst_mult_2_444 ) ) + ( Xd_0__inst_mult_2_302  ) + ( Xd_0__inst_mult_2_301  ))
// Xd_0__inst_mult_2_310  = SHARE((Xd_0__inst_mult_2_440  & Xd_0__inst_mult_2_444 ))

	.dataa(!Xd_0__inst_mult_2_440 ),
	.datab(!Xd_0__inst_mult_2_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_301 ),
	.sharein(Xd_0__inst_mult_2_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_308 ),
	.cout(Xd_0__inst_mult_2_309 ),
	.shareout(Xd_0__inst_mult_2_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_97 (
// Equation(s):
// Xd_0__inst_mult_3_300  = SUM(( !Xd_0__inst_mult_3_428  $ (!Xd_0__inst_mult_3_432  $ (Xd_0__inst_mult_3_39_sumout )) ) + ( Xd_0__inst_mult_3_294  ) + ( Xd_0__inst_mult_3_293  ))
// Xd_0__inst_mult_3_301  = CARRY(( !Xd_0__inst_mult_3_428  $ (!Xd_0__inst_mult_3_432  $ (Xd_0__inst_mult_3_39_sumout )) ) + ( Xd_0__inst_mult_3_294  ) + ( Xd_0__inst_mult_3_293  ))
// Xd_0__inst_mult_3_302  = SHARE((!Xd_0__inst_mult_3_428  & (Xd_0__inst_mult_3_432  & Xd_0__inst_mult_3_39_sumout )) # (Xd_0__inst_mult_3_428  & ((Xd_0__inst_mult_3_39_sumout ) # (Xd_0__inst_mult_3_432 ))))

	.dataa(!Xd_0__inst_mult_3_428 ),
	.datab(!Xd_0__inst_mult_3_432 ),
	.datac(!Xd_0__inst_mult_3_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_293 ),
	.sharein(Xd_0__inst_mult_3_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_300 ),
	.cout(Xd_0__inst_mult_3_301 ),
	.shareout(Xd_0__inst_mult_3_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_98 (
// Equation(s):
// Xd_0__inst_mult_3_304  = SUM(( !Xd_0__inst_mult_3_436  $ (!Xd_0__inst_mult_3_440 ) ) + ( Xd_0__inst_mult_3_298  ) + ( Xd_0__inst_mult_3_297  ))
// Xd_0__inst_mult_3_305  = CARRY(( !Xd_0__inst_mult_3_436  $ (!Xd_0__inst_mult_3_440 ) ) + ( Xd_0__inst_mult_3_298  ) + ( Xd_0__inst_mult_3_297  ))
// Xd_0__inst_mult_3_306  = SHARE((Xd_0__inst_mult_3_436  & Xd_0__inst_mult_3_440 ))

	.dataa(!Xd_0__inst_mult_3_436 ),
	.datab(!Xd_0__inst_mult_3_440 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_297 ),
	.sharein(Xd_0__inst_mult_3_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_304 ),
	.cout(Xd_0__inst_mult_3_305 ),
	.shareout(Xd_0__inst_mult_3_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_101 (
// Equation(s):
// Xd_0__inst_mult_0_304  = SUM(( !Xd_0__inst_mult_0_432  $ (!Xd_0__inst_mult_0_436  $ (Xd_0__inst_mult_0_59_sumout )) ) + ( Xd_0__inst_mult_0_298  ) + ( Xd_0__inst_mult_0_297  ))
// Xd_0__inst_mult_0_305  = CARRY(( !Xd_0__inst_mult_0_432  $ (!Xd_0__inst_mult_0_436  $ (Xd_0__inst_mult_0_59_sumout )) ) + ( Xd_0__inst_mult_0_298  ) + ( Xd_0__inst_mult_0_297  ))
// Xd_0__inst_mult_0_306  = SHARE((!Xd_0__inst_mult_0_432  & (Xd_0__inst_mult_0_436  & Xd_0__inst_mult_0_59_sumout )) # (Xd_0__inst_mult_0_432  & ((Xd_0__inst_mult_0_59_sumout ) # (Xd_0__inst_mult_0_436 ))))

	.dataa(!Xd_0__inst_mult_0_432 ),
	.datab(!Xd_0__inst_mult_0_436 ),
	.datac(!Xd_0__inst_mult_0_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_297 ),
	.sharein(Xd_0__inst_mult_0_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_304 ),
	.cout(Xd_0__inst_mult_0_305 ),
	.shareout(Xd_0__inst_mult_0_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_102 (
// Equation(s):
// Xd_0__inst_mult_0_308  = SUM(( !Xd_0__inst_mult_0_440  $ (!Xd_0__inst_mult_0_444 ) ) + ( Xd_0__inst_mult_0_302  ) + ( Xd_0__inst_mult_0_301  ))
// Xd_0__inst_mult_0_309  = CARRY(( !Xd_0__inst_mult_0_440  $ (!Xd_0__inst_mult_0_444 ) ) + ( Xd_0__inst_mult_0_302  ) + ( Xd_0__inst_mult_0_301  ))
// Xd_0__inst_mult_0_310  = SHARE((Xd_0__inst_mult_0_440  & Xd_0__inst_mult_0_444 ))

	.dataa(!Xd_0__inst_mult_0_440 ),
	.datab(!Xd_0__inst_mult_0_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_301 ),
	.sharein(Xd_0__inst_mult_0_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_308 ),
	.cout(Xd_0__inst_mult_0_309 ),
	.shareout(Xd_0__inst_mult_0_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_101 (
// Equation(s):
// Xd_0__inst_mult_1_304  = SUM(( !Xd_0__inst_mult_1_432  $ (!Xd_0__inst_mult_1_436  $ (Xd_0__inst_mult_1_35_sumout )) ) + ( Xd_0__inst_mult_1_298  ) + ( Xd_0__inst_mult_1_297  ))
// Xd_0__inst_mult_1_305  = CARRY(( !Xd_0__inst_mult_1_432  $ (!Xd_0__inst_mult_1_436  $ (Xd_0__inst_mult_1_35_sumout )) ) + ( Xd_0__inst_mult_1_298  ) + ( Xd_0__inst_mult_1_297  ))
// Xd_0__inst_mult_1_306  = SHARE((!Xd_0__inst_mult_1_432  & (Xd_0__inst_mult_1_436  & Xd_0__inst_mult_1_35_sumout )) # (Xd_0__inst_mult_1_432  & ((Xd_0__inst_mult_1_35_sumout ) # (Xd_0__inst_mult_1_436 ))))

	.dataa(!Xd_0__inst_mult_1_432 ),
	.datab(!Xd_0__inst_mult_1_436 ),
	.datac(!Xd_0__inst_mult_1_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_297 ),
	.sharein(Xd_0__inst_mult_1_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_304 ),
	.cout(Xd_0__inst_mult_1_305 ),
	.shareout(Xd_0__inst_mult_1_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_102 (
// Equation(s):
// Xd_0__inst_mult_1_308  = SUM(( !Xd_0__inst_mult_1_440  $ (!Xd_0__inst_mult_1_444 ) ) + ( Xd_0__inst_mult_1_302  ) + ( Xd_0__inst_mult_1_301  ))
// Xd_0__inst_mult_1_309  = CARRY(( !Xd_0__inst_mult_1_440  $ (!Xd_0__inst_mult_1_444 ) ) + ( Xd_0__inst_mult_1_302  ) + ( Xd_0__inst_mult_1_301  ))
// Xd_0__inst_mult_1_310  = SHARE((Xd_0__inst_mult_1_440  & Xd_0__inst_mult_1_444 ))

	.dataa(!Xd_0__inst_mult_1_440 ),
	.datab(!Xd_0__inst_mult_1_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_301 ),
	.sharein(Xd_0__inst_mult_1_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_308 ),
	.cout(Xd_0__inst_mult_1_309 ),
	.shareout(Xd_0__inst_mult_1_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_111 (
// Equation(s):
// Xd_0__inst_mult_12_356  = SUM(( !Xd_0__inst_mult_12_488  $ (!Xd_0__inst_mult_12_492  $ (Xd_0__inst_mult_12_35_sumout )) ) + ( Xd_0__inst_mult_12_350  ) + ( Xd_0__inst_mult_12_349  ))
// Xd_0__inst_mult_12_357  = CARRY(( !Xd_0__inst_mult_12_488  $ (!Xd_0__inst_mult_12_492  $ (Xd_0__inst_mult_12_35_sumout )) ) + ( Xd_0__inst_mult_12_350  ) + ( Xd_0__inst_mult_12_349  ))
// Xd_0__inst_mult_12_358  = SHARE((!Xd_0__inst_mult_12_488  & (Xd_0__inst_mult_12_492  & Xd_0__inst_mult_12_35_sumout )) # (Xd_0__inst_mult_12_488  & ((Xd_0__inst_mult_12_35_sumout ) # (Xd_0__inst_mult_12_492 ))))

	.dataa(!Xd_0__inst_mult_12_488 ),
	.datab(!Xd_0__inst_mult_12_492 ),
	.datac(!Xd_0__inst_mult_12_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_349 ),
	.sharein(Xd_0__inst_mult_12_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_356 ),
	.cout(Xd_0__inst_mult_12_357 ),
	.shareout(Xd_0__inst_mult_12_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_112 (
// Equation(s):
// Xd_0__inst_mult_12_360  = SUM(( !Xd_0__inst_mult_12_496  $ (!Xd_0__inst_mult_12_500  $ (Xd_0__inst_mult_12_504 )) ) + ( Xd_0__inst_mult_12_354  ) + ( Xd_0__inst_mult_12_353  ))
// Xd_0__inst_mult_12_361  = CARRY(( !Xd_0__inst_mult_12_496  $ (!Xd_0__inst_mult_12_500  $ (Xd_0__inst_mult_12_504 )) ) + ( Xd_0__inst_mult_12_354  ) + ( Xd_0__inst_mult_12_353  ))
// Xd_0__inst_mult_12_362  = SHARE((!Xd_0__inst_mult_12_496  & (Xd_0__inst_mult_12_500  & Xd_0__inst_mult_12_504 )) # (Xd_0__inst_mult_12_496  & ((Xd_0__inst_mult_12_504 ) # (Xd_0__inst_mult_12_500 ))))

	.dataa(!Xd_0__inst_mult_12_496 ),
	.datab(!Xd_0__inst_mult_12_500 ),
	.datac(!Xd_0__inst_mult_12_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_353 ),
	.sharein(Xd_0__inst_mult_12_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_360 ),
	.cout(Xd_0__inst_mult_12_361 ),
	.shareout(Xd_0__inst_mult_12_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_109 (
// Equation(s):
// Xd_0__inst_mult_13_336  = SUM(( !Xd_0__inst_mult_13_464  $ (!Xd_0__inst_mult_13_468  $ (Xd_0__inst_mult_13_39_sumout )) ) + ( Xd_0__inst_mult_13_330  ) + ( Xd_0__inst_mult_13_329  ))
// Xd_0__inst_mult_13_337  = CARRY(( !Xd_0__inst_mult_13_464  $ (!Xd_0__inst_mult_13_468  $ (Xd_0__inst_mult_13_39_sumout )) ) + ( Xd_0__inst_mult_13_330  ) + ( Xd_0__inst_mult_13_329  ))
// Xd_0__inst_mult_13_338  = SHARE((!Xd_0__inst_mult_13_464  & (Xd_0__inst_mult_13_468  & Xd_0__inst_mult_13_39_sumout )) # (Xd_0__inst_mult_13_464  & ((Xd_0__inst_mult_13_39_sumout ) # (Xd_0__inst_mult_13_468 ))))

	.dataa(!Xd_0__inst_mult_13_464 ),
	.datab(!Xd_0__inst_mult_13_468 ),
	.datac(!Xd_0__inst_mult_13_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_329 ),
	.sharein(Xd_0__inst_mult_13_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_336 ),
	.cout(Xd_0__inst_mult_13_337 ),
	.shareout(Xd_0__inst_mult_13_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_110 (
// Equation(s):
// Xd_0__inst_mult_13_340  = SUM(( !Xd_0__inst_mult_13_472  $ (!Xd_0__inst_mult_13_476  $ (Xd_0__inst_mult_13_480 )) ) + ( Xd_0__inst_mult_13_334  ) + ( Xd_0__inst_mult_13_333  ))
// Xd_0__inst_mult_13_341  = CARRY(( !Xd_0__inst_mult_13_472  $ (!Xd_0__inst_mult_13_476  $ (Xd_0__inst_mult_13_480 )) ) + ( Xd_0__inst_mult_13_334  ) + ( Xd_0__inst_mult_13_333  ))
// Xd_0__inst_mult_13_342  = SHARE((!Xd_0__inst_mult_13_472  & (Xd_0__inst_mult_13_476  & Xd_0__inst_mult_13_480 )) # (Xd_0__inst_mult_13_472  & ((Xd_0__inst_mult_13_480 ) # (Xd_0__inst_mult_13_476 ))))

	.dataa(!Xd_0__inst_mult_13_472 ),
	.datab(!Xd_0__inst_mult_13_476 ),
	.datac(!Xd_0__inst_mult_13_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_333 ),
	.sharein(Xd_0__inst_mult_13_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_340 ),
	.cout(Xd_0__inst_mult_13_341 ),
	.shareout(Xd_0__inst_mult_13_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_115 (
// Equation(s):
// Xd_0__inst_mult_14_360  = SUM(( !Xd_0__inst_mult_14_480  $ (!Xd_0__inst_mult_14_484  $ (Xd_0__inst_mult_14_488 )) ) + ( Xd_0__inst_mult_14_358  ) + ( Xd_0__inst_mult_14_357  ))
// Xd_0__inst_mult_14_361  = CARRY(( !Xd_0__inst_mult_14_480  $ (!Xd_0__inst_mult_14_484  $ (Xd_0__inst_mult_14_488 )) ) + ( Xd_0__inst_mult_14_358  ) + ( Xd_0__inst_mult_14_357  ))
// Xd_0__inst_mult_14_362  = SHARE((!Xd_0__inst_mult_14_480  & (Xd_0__inst_mult_14_484  & Xd_0__inst_mult_14_488 )) # (Xd_0__inst_mult_14_480  & ((Xd_0__inst_mult_14_488 ) # (Xd_0__inst_mult_14_484 ))))

	.dataa(!Xd_0__inst_mult_14_480 ),
	.datab(!Xd_0__inst_mult_14_484 ),
	.datac(!Xd_0__inst_mult_14_488 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_357 ),
	.sharein(Xd_0__inst_mult_14_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_360 ),
	.cout(Xd_0__inst_mult_14_361 ),
	.shareout(Xd_0__inst_mult_14_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_115 (
// Equation(s):
// Xd_0__inst_mult_15_360  = SUM(( !Xd_0__inst_mult_15_492  $ (!Xd_0__inst_mult_15_496  $ (Xd_0__inst_mult_15_63_sumout )) ) + ( Xd_0__inst_mult_15_354  ) + ( Xd_0__inst_mult_15_353  ))
// Xd_0__inst_mult_15_361  = CARRY(( !Xd_0__inst_mult_15_492  $ (!Xd_0__inst_mult_15_496  $ (Xd_0__inst_mult_15_63_sumout )) ) + ( Xd_0__inst_mult_15_354  ) + ( Xd_0__inst_mult_15_353  ))
// Xd_0__inst_mult_15_362  = SHARE((!Xd_0__inst_mult_15_492  & (Xd_0__inst_mult_15_496  & Xd_0__inst_mult_15_63_sumout )) # (Xd_0__inst_mult_15_492  & ((Xd_0__inst_mult_15_63_sumout ) # (Xd_0__inst_mult_15_496 ))))

	.dataa(!Xd_0__inst_mult_15_492 ),
	.datab(!Xd_0__inst_mult_15_496 ),
	.datac(!Xd_0__inst_mult_15_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_353 ),
	.sharein(Xd_0__inst_mult_15_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_360 ),
	.cout(Xd_0__inst_mult_15_361 ),
	.shareout(Xd_0__inst_mult_15_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_116 (
// Equation(s):
// Xd_0__inst_mult_15_364  = SUM(( !Xd_0__inst_mult_15_500  $ (!Xd_0__inst_mult_15_504  $ (Xd_0__inst_mult_15_508 )) ) + ( Xd_0__inst_mult_15_358  ) + ( Xd_0__inst_mult_15_357  ))
// Xd_0__inst_mult_15_365  = CARRY(( !Xd_0__inst_mult_15_500  $ (!Xd_0__inst_mult_15_504  $ (Xd_0__inst_mult_15_508 )) ) + ( Xd_0__inst_mult_15_358  ) + ( Xd_0__inst_mult_15_357  ))
// Xd_0__inst_mult_15_366  = SHARE((!Xd_0__inst_mult_15_500  & (Xd_0__inst_mult_15_504  & Xd_0__inst_mult_15_508 )) # (Xd_0__inst_mult_15_500  & ((Xd_0__inst_mult_15_508 ) # (Xd_0__inst_mult_15_504 ))))

	.dataa(!Xd_0__inst_mult_15_500 ),
	.datab(!Xd_0__inst_mult_15_504 ),
	.datac(!Xd_0__inst_mult_15_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_357 ),
	.sharein(Xd_0__inst_mult_15_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_364 ),
	.cout(Xd_0__inst_mult_15_365 ),
	.shareout(Xd_0__inst_mult_15_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_105 (
// Equation(s):
// Xd_0__inst_mult_10_332  = SUM(( !Xd_0__inst_mult_10_460  $ (!Xd_0__inst_mult_10_464  $ (Xd_0__inst_mult_10_59_sumout )) ) + ( Xd_0__inst_mult_10_326  ) + ( Xd_0__inst_mult_10_325  ))
// Xd_0__inst_mult_10_333  = CARRY(( !Xd_0__inst_mult_10_460  $ (!Xd_0__inst_mult_10_464  $ (Xd_0__inst_mult_10_59_sumout )) ) + ( Xd_0__inst_mult_10_326  ) + ( Xd_0__inst_mult_10_325  ))
// Xd_0__inst_mult_10_334  = SHARE((!Xd_0__inst_mult_10_460  & (Xd_0__inst_mult_10_464  & Xd_0__inst_mult_10_59_sumout )) # (Xd_0__inst_mult_10_460  & ((Xd_0__inst_mult_10_59_sumout ) # (Xd_0__inst_mult_10_464 ))))

	.dataa(!Xd_0__inst_mult_10_460 ),
	.datab(!Xd_0__inst_mult_10_464 ),
	.datac(!Xd_0__inst_mult_10_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_325 ),
	.sharein(Xd_0__inst_mult_10_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_332 ),
	.cout(Xd_0__inst_mult_10_333 ),
	.shareout(Xd_0__inst_mult_10_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_106 (
// Equation(s):
// Xd_0__inst_mult_10_336  = SUM(( !Xd_0__inst_mult_10_468  $ (!Xd_0__inst_mult_10_472  $ (Xd_0__inst_mult_10_476 )) ) + ( Xd_0__inst_mult_10_330  ) + ( Xd_0__inst_mult_10_329  ))
// Xd_0__inst_mult_10_337  = CARRY(( !Xd_0__inst_mult_10_468  $ (!Xd_0__inst_mult_10_472  $ (Xd_0__inst_mult_10_476 )) ) + ( Xd_0__inst_mult_10_330  ) + ( Xd_0__inst_mult_10_329  ))
// Xd_0__inst_mult_10_338  = SHARE((!Xd_0__inst_mult_10_468  & (Xd_0__inst_mult_10_472  & Xd_0__inst_mult_10_476 )) # (Xd_0__inst_mult_10_468  & ((Xd_0__inst_mult_10_476 ) # (Xd_0__inst_mult_10_472 ))))

	.dataa(!Xd_0__inst_mult_10_468 ),
	.datab(!Xd_0__inst_mult_10_472 ),
	.datac(!Xd_0__inst_mult_10_476 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_329 ),
	.sharein(Xd_0__inst_mult_10_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_336 ),
	.cout(Xd_0__inst_mult_10_337 ),
	.shareout(Xd_0__inst_mult_10_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_109 (
// Equation(s):
// Xd_0__inst_mult_11_336  = SUM(( !Xd_0__inst_mult_11_464  $ (!Xd_0__inst_mult_11_468  $ (Xd_0__inst_mult_11_55_sumout )) ) + ( Xd_0__inst_mult_11_330  ) + ( Xd_0__inst_mult_11_329  ))
// Xd_0__inst_mult_11_337  = CARRY(( !Xd_0__inst_mult_11_464  $ (!Xd_0__inst_mult_11_468  $ (Xd_0__inst_mult_11_55_sumout )) ) + ( Xd_0__inst_mult_11_330  ) + ( Xd_0__inst_mult_11_329  ))
// Xd_0__inst_mult_11_338  = SHARE((!Xd_0__inst_mult_11_464  & (Xd_0__inst_mult_11_468  & Xd_0__inst_mult_11_55_sumout )) # (Xd_0__inst_mult_11_464  & ((Xd_0__inst_mult_11_55_sumout ) # (Xd_0__inst_mult_11_468 ))))

	.dataa(!Xd_0__inst_mult_11_464 ),
	.datab(!Xd_0__inst_mult_11_468 ),
	.datac(!Xd_0__inst_mult_11_55_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_329 ),
	.sharein(Xd_0__inst_mult_11_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_336 ),
	.cout(Xd_0__inst_mult_11_337 ),
	.shareout(Xd_0__inst_mult_11_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_110 (
// Equation(s):
// Xd_0__inst_mult_11_340  = SUM(( !Xd_0__inst_mult_11_472  $ (!Xd_0__inst_mult_11_476  $ (Xd_0__inst_mult_11_480 )) ) + ( Xd_0__inst_mult_11_334  ) + ( Xd_0__inst_mult_11_333  ))
// Xd_0__inst_mult_11_341  = CARRY(( !Xd_0__inst_mult_11_472  $ (!Xd_0__inst_mult_11_476  $ (Xd_0__inst_mult_11_480 )) ) + ( Xd_0__inst_mult_11_334  ) + ( Xd_0__inst_mult_11_333  ))
// Xd_0__inst_mult_11_342  = SHARE((!Xd_0__inst_mult_11_472  & (Xd_0__inst_mult_11_476  & Xd_0__inst_mult_11_480 )) # (Xd_0__inst_mult_11_472  & ((Xd_0__inst_mult_11_480 ) # (Xd_0__inst_mult_11_476 ))))

	.dataa(!Xd_0__inst_mult_11_472 ),
	.datab(!Xd_0__inst_mult_11_476 ),
	.datac(!Xd_0__inst_mult_11_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_333 ),
	.sharein(Xd_0__inst_mult_11_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_340 ),
	.cout(Xd_0__inst_mult_11_341 ),
	.shareout(Xd_0__inst_mult_11_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_109 (
// Equation(s):
// Xd_0__inst_mult_8_336  = SUM(( !Xd_0__inst_mult_8_464  $ (!Xd_0__inst_mult_8_468  $ (Xd_0__inst_mult_8_35_sumout )) ) + ( Xd_0__inst_mult_8_330  ) + ( Xd_0__inst_mult_8_329  ))
// Xd_0__inst_mult_8_337  = CARRY(( !Xd_0__inst_mult_8_464  $ (!Xd_0__inst_mult_8_468  $ (Xd_0__inst_mult_8_35_sumout )) ) + ( Xd_0__inst_mult_8_330  ) + ( Xd_0__inst_mult_8_329  ))
// Xd_0__inst_mult_8_338  = SHARE((!Xd_0__inst_mult_8_464  & (Xd_0__inst_mult_8_468  & Xd_0__inst_mult_8_35_sumout )) # (Xd_0__inst_mult_8_464  & ((Xd_0__inst_mult_8_35_sumout ) # (Xd_0__inst_mult_8_468 ))))

	.dataa(!Xd_0__inst_mult_8_464 ),
	.datab(!Xd_0__inst_mult_8_468 ),
	.datac(!Xd_0__inst_mult_8_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_329 ),
	.sharein(Xd_0__inst_mult_8_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_336 ),
	.cout(Xd_0__inst_mult_8_337 ),
	.shareout(Xd_0__inst_mult_8_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_110 (
// Equation(s):
// Xd_0__inst_mult_8_340  = SUM(( !Xd_0__inst_mult_8_472  $ (!Xd_0__inst_mult_8_476  $ (Xd_0__inst_mult_8_480 )) ) + ( Xd_0__inst_mult_8_334  ) + ( Xd_0__inst_mult_8_333  ))
// Xd_0__inst_mult_8_341  = CARRY(( !Xd_0__inst_mult_8_472  $ (!Xd_0__inst_mult_8_476  $ (Xd_0__inst_mult_8_480 )) ) + ( Xd_0__inst_mult_8_334  ) + ( Xd_0__inst_mult_8_333  ))
// Xd_0__inst_mult_8_342  = SHARE((!Xd_0__inst_mult_8_472  & (Xd_0__inst_mult_8_476  & Xd_0__inst_mult_8_480 )) # (Xd_0__inst_mult_8_472  & ((Xd_0__inst_mult_8_480 ) # (Xd_0__inst_mult_8_476 ))))

	.dataa(!Xd_0__inst_mult_8_472 ),
	.datab(!Xd_0__inst_mult_8_476 ),
	.datac(!Xd_0__inst_mult_8_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_333 ),
	.sharein(Xd_0__inst_mult_8_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_340 ),
	.cout(Xd_0__inst_mult_8_341 ),
	.shareout(Xd_0__inst_mult_8_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_105 (
// Equation(s):
// Xd_0__inst_mult_9_332  = SUM(( !Xd_0__inst_mult_9_460  $ (!Xd_0__inst_mult_9_464  $ (Xd_0__inst_mult_9_55_sumout )) ) + ( Xd_0__inst_mult_9_326  ) + ( Xd_0__inst_mult_9_325  ))
// Xd_0__inst_mult_9_333  = CARRY(( !Xd_0__inst_mult_9_460  $ (!Xd_0__inst_mult_9_464  $ (Xd_0__inst_mult_9_55_sumout )) ) + ( Xd_0__inst_mult_9_326  ) + ( Xd_0__inst_mult_9_325  ))
// Xd_0__inst_mult_9_334  = SHARE((!Xd_0__inst_mult_9_460  & (Xd_0__inst_mult_9_464  & Xd_0__inst_mult_9_55_sumout )) # (Xd_0__inst_mult_9_460  & ((Xd_0__inst_mult_9_55_sumout ) # (Xd_0__inst_mult_9_464 ))))

	.dataa(!Xd_0__inst_mult_9_460 ),
	.datab(!Xd_0__inst_mult_9_464 ),
	.datac(!Xd_0__inst_mult_9_55_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_325 ),
	.sharein(Xd_0__inst_mult_9_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_332 ),
	.cout(Xd_0__inst_mult_9_333 ),
	.shareout(Xd_0__inst_mult_9_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_106 (
// Equation(s):
// Xd_0__inst_mult_9_336  = SUM(( !Xd_0__inst_mult_9_468  $ (!Xd_0__inst_mult_9_472  $ (Xd_0__inst_mult_9_476 )) ) + ( Xd_0__inst_mult_9_330  ) + ( Xd_0__inst_mult_9_329  ))
// Xd_0__inst_mult_9_337  = CARRY(( !Xd_0__inst_mult_9_468  $ (!Xd_0__inst_mult_9_472  $ (Xd_0__inst_mult_9_476 )) ) + ( Xd_0__inst_mult_9_330  ) + ( Xd_0__inst_mult_9_329  ))
// Xd_0__inst_mult_9_338  = SHARE((!Xd_0__inst_mult_9_468  & (Xd_0__inst_mult_9_472  & Xd_0__inst_mult_9_476 )) # (Xd_0__inst_mult_9_468  & ((Xd_0__inst_mult_9_476 ) # (Xd_0__inst_mult_9_472 ))))

	.dataa(!Xd_0__inst_mult_9_468 ),
	.datab(!Xd_0__inst_mult_9_472 ),
	.datac(!Xd_0__inst_mult_9_476 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_329 ),
	.sharein(Xd_0__inst_mult_9_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_336 ),
	.cout(Xd_0__inst_mult_9_337 ),
	.shareout(Xd_0__inst_mult_9_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_105 (
// Equation(s):
// Xd_0__inst_mult_6_332  = SUM(( !Xd_0__inst_mult_6_460  $ (!Xd_0__inst_mult_6_464  $ (Xd_0__inst_mult_6_35_sumout )) ) + ( Xd_0__inst_mult_6_326  ) + ( Xd_0__inst_mult_6_325  ))
// Xd_0__inst_mult_6_333  = CARRY(( !Xd_0__inst_mult_6_460  $ (!Xd_0__inst_mult_6_464  $ (Xd_0__inst_mult_6_35_sumout )) ) + ( Xd_0__inst_mult_6_326  ) + ( Xd_0__inst_mult_6_325  ))
// Xd_0__inst_mult_6_334  = SHARE((!Xd_0__inst_mult_6_460  & (Xd_0__inst_mult_6_464  & Xd_0__inst_mult_6_35_sumout )) # (Xd_0__inst_mult_6_460  & ((Xd_0__inst_mult_6_35_sumout ) # (Xd_0__inst_mult_6_464 ))))

	.dataa(!Xd_0__inst_mult_6_460 ),
	.datab(!Xd_0__inst_mult_6_464 ),
	.datac(!Xd_0__inst_mult_6_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_325 ),
	.sharein(Xd_0__inst_mult_6_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_332 ),
	.cout(Xd_0__inst_mult_6_333 ),
	.shareout(Xd_0__inst_mult_6_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_106 (
// Equation(s):
// Xd_0__inst_mult_6_336  = SUM(( !Xd_0__inst_mult_6_468  $ (!Xd_0__inst_mult_6_472  $ (Xd_0__inst_mult_6_476 )) ) + ( Xd_0__inst_mult_6_330  ) + ( Xd_0__inst_mult_6_329  ))
// Xd_0__inst_mult_6_337  = CARRY(( !Xd_0__inst_mult_6_468  $ (!Xd_0__inst_mult_6_472  $ (Xd_0__inst_mult_6_476 )) ) + ( Xd_0__inst_mult_6_330  ) + ( Xd_0__inst_mult_6_329  ))
// Xd_0__inst_mult_6_338  = SHARE((!Xd_0__inst_mult_6_468  & (Xd_0__inst_mult_6_472  & Xd_0__inst_mult_6_476 )) # (Xd_0__inst_mult_6_468  & ((Xd_0__inst_mult_6_476 ) # (Xd_0__inst_mult_6_472 ))))

	.dataa(!Xd_0__inst_mult_6_468 ),
	.datab(!Xd_0__inst_mult_6_472 ),
	.datac(!Xd_0__inst_mult_6_476 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_329 ),
	.sharein(Xd_0__inst_mult_6_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_336 ),
	.cout(Xd_0__inst_mult_6_337 ),
	.shareout(Xd_0__inst_mult_6_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_99 (
// Equation(s):
// Xd_0__inst_mult_7_308  = SUM(( !Xd_0__inst_mult_7_444  $ (!Xd_0__inst_mult_7_448  $ (Xd_0__inst_mult_7_35_sumout )) ) + ( Xd_0__inst_mult_7_302  ) + ( Xd_0__inst_mult_7_301  ))
// Xd_0__inst_mult_7_309  = CARRY(( !Xd_0__inst_mult_7_444  $ (!Xd_0__inst_mult_7_448  $ (Xd_0__inst_mult_7_35_sumout )) ) + ( Xd_0__inst_mult_7_302  ) + ( Xd_0__inst_mult_7_301  ))
// Xd_0__inst_mult_7_310  = SHARE((!Xd_0__inst_mult_7_444  & (Xd_0__inst_mult_7_448  & Xd_0__inst_mult_7_35_sumout )) # (Xd_0__inst_mult_7_444  & ((Xd_0__inst_mult_7_35_sumout ) # (Xd_0__inst_mult_7_448 ))))

	.dataa(!Xd_0__inst_mult_7_444 ),
	.datab(!Xd_0__inst_mult_7_448 ),
	.datac(!Xd_0__inst_mult_7_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_301 ),
	.sharein(Xd_0__inst_mult_7_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_308 ),
	.cout(Xd_0__inst_mult_7_309 ),
	.shareout(Xd_0__inst_mult_7_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_100 (
// Equation(s):
// Xd_0__inst_mult_7_312  = SUM(( !Xd_0__inst_mult_7_452  $ (!Xd_0__inst_mult_7_456  $ (Xd_0__inst_mult_7_460 )) ) + ( Xd_0__inst_mult_7_306  ) + ( Xd_0__inst_mult_7_305  ))
// Xd_0__inst_mult_7_313  = CARRY(( !Xd_0__inst_mult_7_452  $ (!Xd_0__inst_mult_7_456  $ (Xd_0__inst_mult_7_460 )) ) + ( Xd_0__inst_mult_7_306  ) + ( Xd_0__inst_mult_7_305  ))
// Xd_0__inst_mult_7_314  = SHARE((!Xd_0__inst_mult_7_452  & (Xd_0__inst_mult_7_456  & Xd_0__inst_mult_7_460 )) # (Xd_0__inst_mult_7_452  & ((Xd_0__inst_mult_7_460 ) # (Xd_0__inst_mult_7_456 ))))

	.dataa(!Xd_0__inst_mult_7_452 ),
	.datab(!Xd_0__inst_mult_7_456 ),
	.datac(!Xd_0__inst_mult_7_460 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_305 ),
	.sharein(Xd_0__inst_mult_7_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_312 ),
	.cout(Xd_0__inst_mult_7_313 ),
	.shareout(Xd_0__inst_mult_7_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_111 (
// Equation(s):
// Xd_0__inst_mult_4_344  = SUM(( !Xd_0__inst_mult_4_484  $ (!Xd_0__inst_mult_4_488  $ (Xd_0__inst_mult_4_55_sumout )) ) + ( Xd_0__inst_mult_4_338  ) + ( Xd_0__inst_mult_4_337  ))
// Xd_0__inst_mult_4_345  = CARRY(( !Xd_0__inst_mult_4_484  $ (!Xd_0__inst_mult_4_488  $ (Xd_0__inst_mult_4_55_sumout )) ) + ( Xd_0__inst_mult_4_338  ) + ( Xd_0__inst_mult_4_337  ))
// Xd_0__inst_mult_4_346  = SHARE((!Xd_0__inst_mult_4_484  & (Xd_0__inst_mult_4_488  & Xd_0__inst_mult_4_55_sumout )) # (Xd_0__inst_mult_4_484  & ((Xd_0__inst_mult_4_55_sumout ) # (Xd_0__inst_mult_4_488 ))))

	.dataa(!Xd_0__inst_mult_4_484 ),
	.datab(!Xd_0__inst_mult_4_488 ),
	.datac(!Xd_0__inst_mult_4_55_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_337 ),
	.sharein(Xd_0__inst_mult_4_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_344 ),
	.cout(Xd_0__inst_mult_4_345 ),
	.shareout(Xd_0__inst_mult_4_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_112 (
// Equation(s):
// Xd_0__inst_mult_4_348  = SUM(( !Xd_0__inst_mult_4_492  $ (!Xd_0__inst_mult_4_496  $ (Xd_0__inst_mult_4_500 )) ) + ( Xd_0__inst_mult_4_342  ) + ( Xd_0__inst_mult_4_341  ))
// Xd_0__inst_mult_4_349  = CARRY(( !Xd_0__inst_mult_4_492  $ (!Xd_0__inst_mult_4_496  $ (Xd_0__inst_mult_4_500 )) ) + ( Xd_0__inst_mult_4_342  ) + ( Xd_0__inst_mult_4_341  ))
// Xd_0__inst_mult_4_350  = SHARE((!Xd_0__inst_mult_4_492  & (Xd_0__inst_mult_4_496  & Xd_0__inst_mult_4_500 )) # (Xd_0__inst_mult_4_492  & ((Xd_0__inst_mult_4_500 ) # (Xd_0__inst_mult_4_496 ))))

	.dataa(!Xd_0__inst_mult_4_492 ),
	.datab(!Xd_0__inst_mult_4_496 ),
	.datac(!Xd_0__inst_mult_4_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_341 ),
	.sharein(Xd_0__inst_mult_4_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_348 ),
	.cout(Xd_0__inst_mult_4_349 ),
	.shareout(Xd_0__inst_mult_4_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_99 (
// Equation(s):
// Xd_0__inst_mult_5_308  = SUM(( !Xd_0__inst_mult_5_444  $ (!Xd_0__inst_mult_5_448  $ (Xd_0__inst_mult_7_380 )) ) + ( Xd_0__inst_mult_5_302  ) + ( Xd_0__inst_mult_5_301  ))
// Xd_0__inst_mult_5_309  = CARRY(( !Xd_0__inst_mult_5_444  $ (!Xd_0__inst_mult_5_448  $ (Xd_0__inst_mult_7_380 )) ) + ( Xd_0__inst_mult_5_302  ) + ( Xd_0__inst_mult_5_301  ))
// Xd_0__inst_mult_5_310  = SHARE((!Xd_0__inst_mult_5_444  & (Xd_0__inst_mult_5_448  & Xd_0__inst_mult_7_380 )) # (Xd_0__inst_mult_5_444  & ((Xd_0__inst_mult_7_380 ) # (Xd_0__inst_mult_5_448 ))))

	.dataa(!Xd_0__inst_mult_5_444 ),
	.datab(!Xd_0__inst_mult_5_448 ),
	.datac(!Xd_0__inst_mult_7_380 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_301 ),
	.sharein(Xd_0__inst_mult_5_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_308 ),
	.cout(Xd_0__inst_mult_5_309 ),
	.shareout(Xd_0__inst_mult_5_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_100 (
// Equation(s):
// Xd_0__inst_mult_5_312  = SUM(( !Xd_0__inst_mult_5_452  $ (!Xd_0__inst_mult_5_456  $ (Xd_0__inst_mult_5_460 )) ) + ( Xd_0__inst_mult_5_306  ) + ( Xd_0__inst_mult_5_305  ))
// Xd_0__inst_mult_5_313  = CARRY(( !Xd_0__inst_mult_5_452  $ (!Xd_0__inst_mult_5_456  $ (Xd_0__inst_mult_5_460 )) ) + ( Xd_0__inst_mult_5_306  ) + ( Xd_0__inst_mult_5_305  ))
// Xd_0__inst_mult_5_314  = SHARE((!Xd_0__inst_mult_5_452  & (Xd_0__inst_mult_5_456  & Xd_0__inst_mult_5_460 )) # (Xd_0__inst_mult_5_452  & ((Xd_0__inst_mult_5_460 ) # (Xd_0__inst_mult_5_456 ))))

	.dataa(!Xd_0__inst_mult_5_452 ),
	.datab(!Xd_0__inst_mult_5_456 ),
	.datac(!Xd_0__inst_mult_5_460 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_305 ),
	.sharein(Xd_0__inst_mult_5_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_312 ),
	.cout(Xd_0__inst_mult_5_313 ),
	.shareout(Xd_0__inst_mult_5_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_103 (
// Equation(s):
// Xd_0__inst_mult_2_312  = SUM(( !Xd_0__inst_mult_2_448  $ (!Xd_0__inst_mult_2_452  $ (Xd_0__inst_mult_2_67_sumout )) ) + ( Xd_0__inst_mult_2_306  ) + ( Xd_0__inst_mult_2_305  ))
// Xd_0__inst_mult_2_313  = CARRY(( !Xd_0__inst_mult_2_448  $ (!Xd_0__inst_mult_2_452  $ (Xd_0__inst_mult_2_67_sumout )) ) + ( Xd_0__inst_mult_2_306  ) + ( Xd_0__inst_mult_2_305  ))
// Xd_0__inst_mult_2_314  = SHARE((!Xd_0__inst_mult_2_448  & (Xd_0__inst_mult_2_452  & Xd_0__inst_mult_2_67_sumout )) # (Xd_0__inst_mult_2_448  & ((Xd_0__inst_mult_2_67_sumout ) # (Xd_0__inst_mult_2_452 ))))

	.dataa(!Xd_0__inst_mult_2_448 ),
	.datab(!Xd_0__inst_mult_2_452 ),
	.datac(!Xd_0__inst_mult_2_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_305 ),
	.sharein(Xd_0__inst_mult_2_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_312 ),
	.cout(Xd_0__inst_mult_2_313 ),
	.shareout(Xd_0__inst_mult_2_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_104 (
// Equation(s):
// Xd_0__inst_mult_2_316  = SUM(( !Xd_0__inst_mult_2_456  $ (!Xd_0__inst_mult_2_460  $ (Xd_0__inst_mult_2_464 )) ) + ( Xd_0__inst_mult_2_310  ) + ( Xd_0__inst_mult_2_309  ))
// Xd_0__inst_mult_2_317  = CARRY(( !Xd_0__inst_mult_2_456  $ (!Xd_0__inst_mult_2_460  $ (Xd_0__inst_mult_2_464 )) ) + ( Xd_0__inst_mult_2_310  ) + ( Xd_0__inst_mult_2_309  ))
// Xd_0__inst_mult_2_318  = SHARE((!Xd_0__inst_mult_2_456  & (Xd_0__inst_mult_2_460  & Xd_0__inst_mult_2_464 )) # (Xd_0__inst_mult_2_456  & ((Xd_0__inst_mult_2_464 ) # (Xd_0__inst_mult_2_460 ))))

	.dataa(!Xd_0__inst_mult_2_456 ),
	.datab(!Xd_0__inst_mult_2_460 ),
	.datac(!Xd_0__inst_mult_2_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_309 ),
	.sharein(Xd_0__inst_mult_2_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_316 ),
	.cout(Xd_0__inst_mult_2_317 ),
	.shareout(Xd_0__inst_mult_2_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_99 (
// Equation(s):
// Xd_0__inst_mult_3_308  = SUM(( !Xd_0__inst_mult_3_444  $ (!Xd_0__inst_mult_3_448  $ (Xd_0__inst_mult_3_63_sumout )) ) + ( Xd_0__inst_mult_3_302  ) + ( Xd_0__inst_mult_3_301  ))
// Xd_0__inst_mult_3_309  = CARRY(( !Xd_0__inst_mult_3_444  $ (!Xd_0__inst_mult_3_448  $ (Xd_0__inst_mult_3_63_sumout )) ) + ( Xd_0__inst_mult_3_302  ) + ( Xd_0__inst_mult_3_301  ))
// Xd_0__inst_mult_3_310  = SHARE((!Xd_0__inst_mult_3_444  & (Xd_0__inst_mult_3_448  & Xd_0__inst_mult_3_63_sumout )) # (Xd_0__inst_mult_3_444  & ((Xd_0__inst_mult_3_63_sumout ) # (Xd_0__inst_mult_3_448 ))))

	.dataa(!Xd_0__inst_mult_3_444 ),
	.datab(!Xd_0__inst_mult_3_448 ),
	.datac(!Xd_0__inst_mult_3_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_301 ),
	.sharein(Xd_0__inst_mult_3_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_308 ),
	.cout(Xd_0__inst_mult_3_309 ),
	.shareout(Xd_0__inst_mult_3_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_100 (
// Equation(s):
// Xd_0__inst_mult_3_312  = SUM(( !Xd_0__inst_mult_3_452  $ (!Xd_0__inst_mult_3_456  $ (Xd_0__inst_mult_3_460 )) ) + ( Xd_0__inst_mult_3_306  ) + ( Xd_0__inst_mult_3_305  ))
// Xd_0__inst_mult_3_313  = CARRY(( !Xd_0__inst_mult_3_452  $ (!Xd_0__inst_mult_3_456  $ (Xd_0__inst_mult_3_460 )) ) + ( Xd_0__inst_mult_3_306  ) + ( Xd_0__inst_mult_3_305  ))
// Xd_0__inst_mult_3_314  = SHARE((!Xd_0__inst_mult_3_452  & (Xd_0__inst_mult_3_456  & Xd_0__inst_mult_3_460 )) # (Xd_0__inst_mult_3_452  & ((Xd_0__inst_mult_3_460 ) # (Xd_0__inst_mult_3_456 ))))

	.dataa(!Xd_0__inst_mult_3_452 ),
	.datab(!Xd_0__inst_mult_3_456 ),
	.datac(!Xd_0__inst_mult_3_460 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_305 ),
	.sharein(Xd_0__inst_mult_3_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_312 ),
	.cout(Xd_0__inst_mult_3_313 ),
	.shareout(Xd_0__inst_mult_3_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_103 (
// Equation(s):
// Xd_0__inst_mult_0_312  = SUM(( !Xd_0__inst_mult_0_448  $ (!Xd_0__inst_mult_0_452  $ (Xd_0__inst_mult_0_67_sumout )) ) + ( Xd_0__inst_mult_0_306  ) + ( Xd_0__inst_mult_0_305  ))
// Xd_0__inst_mult_0_313  = CARRY(( !Xd_0__inst_mult_0_448  $ (!Xd_0__inst_mult_0_452  $ (Xd_0__inst_mult_0_67_sumout )) ) + ( Xd_0__inst_mult_0_306  ) + ( Xd_0__inst_mult_0_305  ))
// Xd_0__inst_mult_0_314  = SHARE((!Xd_0__inst_mult_0_448  & (Xd_0__inst_mult_0_452  & Xd_0__inst_mult_0_67_sumout )) # (Xd_0__inst_mult_0_448  & ((Xd_0__inst_mult_0_67_sumout ) # (Xd_0__inst_mult_0_452 ))))

	.dataa(!Xd_0__inst_mult_0_448 ),
	.datab(!Xd_0__inst_mult_0_452 ),
	.datac(!Xd_0__inst_mult_0_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_305 ),
	.sharein(Xd_0__inst_mult_0_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_312 ),
	.cout(Xd_0__inst_mult_0_313 ),
	.shareout(Xd_0__inst_mult_0_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_104 (
// Equation(s):
// Xd_0__inst_mult_0_316  = SUM(( !Xd_0__inst_mult_0_456  $ (!Xd_0__inst_mult_0_460  $ (Xd_0__inst_mult_0_464 )) ) + ( Xd_0__inst_mult_0_310  ) + ( Xd_0__inst_mult_0_309  ))
// Xd_0__inst_mult_0_317  = CARRY(( !Xd_0__inst_mult_0_456  $ (!Xd_0__inst_mult_0_460  $ (Xd_0__inst_mult_0_464 )) ) + ( Xd_0__inst_mult_0_310  ) + ( Xd_0__inst_mult_0_309  ))
// Xd_0__inst_mult_0_318  = SHARE((!Xd_0__inst_mult_0_456  & (Xd_0__inst_mult_0_460  & Xd_0__inst_mult_0_464 )) # (Xd_0__inst_mult_0_456  & ((Xd_0__inst_mult_0_464 ) # (Xd_0__inst_mult_0_460 ))))

	.dataa(!Xd_0__inst_mult_0_456 ),
	.datab(!Xd_0__inst_mult_0_460 ),
	.datac(!Xd_0__inst_mult_0_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_309 ),
	.sharein(Xd_0__inst_mult_0_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_316 ),
	.cout(Xd_0__inst_mult_0_317 ),
	.shareout(Xd_0__inst_mult_0_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_103 (
// Equation(s):
// Xd_0__inst_mult_1_312  = SUM(( !Xd_0__inst_mult_1_448  $ (!Xd_0__inst_mult_1_452  $ (Xd_0__inst_mult_1_39_sumout )) ) + ( Xd_0__inst_mult_1_306  ) + ( Xd_0__inst_mult_1_305  ))
// Xd_0__inst_mult_1_313  = CARRY(( !Xd_0__inst_mult_1_448  $ (!Xd_0__inst_mult_1_452  $ (Xd_0__inst_mult_1_39_sumout )) ) + ( Xd_0__inst_mult_1_306  ) + ( Xd_0__inst_mult_1_305  ))
// Xd_0__inst_mult_1_314  = SHARE((!Xd_0__inst_mult_1_448  & (Xd_0__inst_mult_1_452  & Xd_0__inst_mult_1_39_sumout )) # (Xd_0__inst_mult_1_448  & ((Xd_0__inst_mult_1_39_sumout ) # (Xd_0__inst_mult_1_452 ))))

	.dataa(!Xd_0__inst_mult_1_448 ),
	.datab(!Xd_0__inst_mult_1_452 ),
	.datac(!Xd_0__inst_mult_1_39_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_305 ),
	.sharein(Xd_0__inst_mult_1_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_312 ),
	.cout(Xd_0__inst_mult_1_313 ),
	.shareout(Xd_0__inst_mult_1_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_104 (
// Equation(s):
// Xd_0__inst_mult_1_316  = SUM(( !Xd_0__inst_mult_1_456  $ (!Xd_0__inst_mult_1_460  $ (Xd_0__inst_mult_1_464 )) ) + ( Xd_0__inst_mult_1_310  ) + ( Xd_0__inst_mult_1_309  ))
// Xd_0__inst_mult_1_317  = CARRY(( !Xd_0__inst_mult_1_456  $ (!Xd_0__inst_mult_1_460  $ (Xd_0__inst_mult_1_464 )) ) + ( Xd_0__inst_mult_1_310  ) + ( Xd_0__inst_mult_1_309  ))
// Xd_0__inst_mult_1_318  = SHARE((!Xd_0__inst_mult_1_456  & (Xd_0__inst_mult_1_460  & Xd_0__inst_mult_1_464 )) # (Xd_0__inst_mult_1_456  & ((Xd_0__inst_mult_1_464 ) # (Xd_0__inst_mult_1_460 ))))

	.dataa(!Xd_0__inst_mult_1_456 ),
	.datab(!Xd_0__inst_mult_1_460 ),
	.datac(!Xd_0__inst_mult_1_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_309 ),
	.sharein(Xd_0__inst_mult_1_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_316 ),
	.cout(Xd_0__inst_mult_1_317 ),
	.shareout(Xd_0__inst_mult_1_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_113 (
// Equation(s):
// Xd_0__inst_mult_12_364  = SUM(( !Xd_0__inst_mult_12_508  $ (!Xd_0__inst_mult_12_512 ) ) + ( Xd_0__inst_mult_12_358  ) + ( Xd_0__inst_mult_12_357  ))
// Xd_0__inst_mult_12_365  = CARRY(( !Xd_0__inst_mult_12_508  $ (!Xd_0__inst_mult_12_512 ) ) + ( Xd_0__inst_mult_12_358  ) + ( Xd_0__inst_mult_12_357  ))
// Xd_0__inst_mult_12_366  = SHARE((Xd_0__inst_mult_12_508  & Xd_0__inst_mult_12_512 ))

	.dataa(!Xd_0__inst_mult_12_508 ),
	.datab(!Xd_0__inst_mult_12_512 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_357 ),
	.sharein(Xd_0__inst_mult_12_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_364 ),
	.cout(Xd_0__inst_mult_12_365 ),
	.shareout(Xd_0__inst_mult_12_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_114 (
// Equation(s):
// Xd_0__inst_mult_12_368  = SUM(( !Xd_0__inst_mult_12_516  $ (!Xd_0__inst_mult_12_520  $ (Xd_0__inst_mult_12_524 )) ) + ( Xd_0__inst_mult_12_362  ) + ( Xd_0__inst_mult_12_361  ))
// Xd_0__inst_mult_12_369  = CARRY(( !Xd_0__inst_mult_12_516  $ (!Xd_0__inst_mult_12_520  $ (Xd_0__inst_mult_12_524 )) ) + ( Xd_0__inst_mult_12_362  ) + ( Xd_0__inst_mult_12_361  ))
// Xd_0__inst_mult_12_370  = SHARE((!Xd_0__inst_mult_12_516  & (Xd_0__inst_mult_12_520  & Xd_0__inst_mult_12_524 )) # (Xd_0__inst_mult_12_516  & ((Xd_0__inst_mult_12_524 ) # (Xd_0__inst_mult_12_520 ))))

	.dataa(!Xd_0__inst_mult_12_516 ),
	.datab(!Xd_0__inst_mult_12_520 ),
	.datac(!Xd_0__inst_mult_12_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_361 ),
	.sharein(Xd_0__inst_mult_12_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_368 ),
	.cout(Xd_0__inst_mult_12_369 ),
	.shareout(Xd_0__inst_mult_12_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_111 (
// Equation(s):
// Xd_0__inst_mult_13_344  = SUM(( !Xd_0__inst_mult_13_484  $ (!Xd_0__inst_mult_13_488 ) ) + ( Xd_0__inst_mult_13_338  ) + ( Xd_0__inst_mult_13_337  ))
// Xd_0__inst_mult_13_345  = CARRY(( !Xd_0__inst_mult_13_484  $ (!Xd_0__inst_mult_13_488 ) ) + ( Xd_0__inst_mult_13_338  ) + ( Xd_0__inst_mult_13_337  ))
// Xd_0__inst_mult_13_346  = SHARE((Xd_0__inst_mult_13_484  & Xd_0__inst_mult_13_488 ))

	.dataa(!Xd_0__inst_mult_13_484 ),
	.datab(!Xd_0__inst_mult_13_488 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_337 ),
	.sharein(Xd_0__inst_mult_13_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_344 ),
	.cout(Xd_0__inst_mult_13_345 ),
	.shareout(Xd_0__inst_mult_13_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_112 (
// Equation(s):
// Xd_0__inst_mult_13_348  = SUM(( !Xd_0__inst_mult_13_492  $ (!Xd_0__inst_mult_13_496  $ (Xd_0__inst_mult_13_500 )) ) + ( Xd_0__inst_mult_13_342  ) + ( Xd_0__inst_mult_13_341  ))
// Xd_0__inst_mult_13_349  = CARRY(( !Xd_0__inst_mult_13_492  $ (!Xd_0__inst_mult_13_496  $ (Xd_0__inst_mult_13_500 )) ) + ( Xd_0__inst_mult_13_342  ) + ( Xd_0__inst_mult_13_341  ))
// Xd_0__inst_mult_13_350  = SHARE((!Xd_0__inst_mult_13_492  & (Xd_0__inst_mult_13_496  & Xd_0__inst_mult_13_500 )) # (Xd_0__inst_mult_13_492  & ((Xd_0__inst_mult_13_500 ) # (Xd_0__inst_mult_13_496 ))))

	.dataa(!Xd_0__inst_mult_13_492 ),
	.datab(!Xd_0__inst_mult_13_496 ),
	.datac(!Xd_0__inst_mult_13_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_341 ),
	.sharein(Xd_0__inst_mult_13_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_348 ),
	.cout(Xd_0__inst_mult_13_349 ),
	.shareout(Xd_0__inst_mult_13_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_116 (
// Equation(s):
// Xd_0__inst_mult_14_364  = SUM(( !Xd_0__inst_mult_14_492  $ (!Xd_0__inst_mult_14_496  $ (Xd_0__inst_mult_14_500 )) ) + ( Xd_0__inst_mult_14_362  ) + ( Xd_0__inst_mult_14_361  ))
// Xd_0__inst_mult_14_365  = CARRY(( !Xd_0__inst_mult_14_492  $ (!Xd_0__inst_mult_14_496  $ (Xd_0__inst_mult_14_500 )) ) + ( Xd_0__inst_mult_14_362  ) + ( Xd_0__inst_mult_14_361  ))
// Xd_0__inst_mult_14_366  = SHARE((!Xd_0__inst_mult_14_492  & (Xd_0__inst_mult_14_496  & Xd_0__inst_mult_14_500 )) # (Xd_0__inst_mult_14_492  & ((Xd_0__inst_mult_14_500 ) # (Xd_0__inst_mult_14_496 ))))

	.dataa(!Xd_0__inst_mult_14_492 ),
	.datab(!Xd_0__inst_mult_14_496 ),
	.datac(!Xd_0__inst_mult_14_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_361 ),
	.sharein(Xd_0__inst_mult_14_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_364 ),
	.cout(Xd_0__inst_mult_14_365 ),
	.shareout(Xd_0__inst_mult_14_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_117 (
// Equation(s):
// Xd_0__inst_mult_15_368  = SUM(( !Xd_0__inst_mult_15_512  $ (!Xd_0__inst_mult_15_516 ) ) + ( Xd_0__inst_mult_15_362  ) + ( Xd_0__inst_mult_15_361  ))
// Xd_0__inst_mult_15_369  = CARRY(( !Xd_0__inst_mult_15_512  $ (!Xd_0__inst_mult_15_516 ) ) + ( Xd_0__inst_mult_15_362  ) + ( Xd_0__inst_mult_15_361  ))
// Xd_0__inst_mult_15_370  = SHARE((Xd_0__inst_mult_15_512  & Xd_0__inst_mult_15_516 ))

	.dataa(!Xd_0__inst_mult_15_512 ),
	.datab(!Xd_0__inst_mult_15_516 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_361 ),
	.sharein(Xd_0__inst_mult_15_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_368 ),
	.cout(Xd_0__inst_mult_15_369 ),
	.shareout(Xd_0__inst_mult_15_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_118 (
// Equation(s):
// Xd_0__inst_mult_15_372  = SUM(( !Xd_0__inst_mult_15_520  $ (!Xd_0__inst_mult_15_524  $ (Xd_0__inst_mult_15_528 )) ) + ( Xd_0__inst_mult_15_366  ) + ( Xd_0__inst_mult_15_365  ))
// Xd_0__inst_mult_15_373  = CARRY(( !Xd_0__inst_mult_15_520  $ (!Xd_0__inst_mult_15_524  $ (Xd_0__inst_mult_15_528 )) ) + ( Xd_0__inst_mult_15_366  ) + ( Xd_0__inst_mult_15_365  ))
// Xd_0__inst_mult_15_374  = SHARE((!Xd_0__inst_mult_15_520  & (Xd_0__inst_mult_15_524  & Xd_0__inst_mult_15_528 )) # (Xd_0__inst_mult_15_520  & ((Xd_0__inst_mult_15_528 ) # (Xd_0__inst_mult_15_524 ))))

	.dataa(!Xd_0__inst_mult_15_520 ),
	.datab(!Xd_0__inst_mult_15_524 ),
	.datac(!Xd_0__inst_mult_15_528 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_365 ),
	.sharein(Xd_0__inst_mult_15_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_372 ),
	.cout(Xd_0__inst_mult_15_373 ),
	.shareout(Xd_0__inst_mult_15_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_107 (
// Equation(s):
// Xd_0__inst_mult_10_340  = SUM(( !Xd_0__inst_mult_10_480  $ (!Xd_0__inst_mult_10_484 ) ) + ( Xd_0__inst_mult_10_334  ) + ( Xd_0__inst_mult_10_333  ))
// Xd_0__inst_mult_10_341  = CARRY(( !Xd_0__inst_mult_10_480  $ (!Xd_0__inst_mult_10_484 ) ) + ( Xd_0__inst_mult_10_334  ) + ( Xd_0__inst_mult_10_333  ))
// Xd_0__inst_mult_10_342  = SHARE((Xd_0__inst_mult_10_480  & Xd_0__inst_mult_10_484 ))

	.dataa(!Xd_0__inst_mult_10_480 ),
	.datab(!Xd_0__inst_mult_10_484 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_333 ),
	.sharein(Xd_0__inst_mult_10_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_340 ),
	.cout(Xd_0__inst_mult_10_341 ),
	.shareout(Xd_0__inst_mult_10_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_108 (
// Equation(s):
// Xd_0__inst_mult_10_344  = SUM(( !Xd_0__inst_mult_10_488  $ (!Xd_0__inst_mult_10_492  $ (Xd_0__inst_mult_10_496 )) ) + ( Xd_0__inst_mult_10_338  ) + ( Xd_0__inst_mult_10_337  ))
// Xd_0__inst_mult_10_345  = CARRY(( !Xd_0__inst_mult_10_488  $ (!Xd_0__inst_mult_10_492  $ (Xd_0__inst_mult_10_496 )) ) + ( Xd_0__inst_mult_10_338  ) + ( Xd_0__inst_mult_10_337  ))
// Xd_0__inst_mult_10_346  = SHARE((!Xd_0__inst_mult_10_488  & (Xd_0__inst_mult_10_492  & Xd_0__inst_mult_10_496 )) # (Xd_0__inst_mult_10_488  & ((Xd_0__inst_mult_10_496 ) # (Xd_0__inst_mult_10_492 ))))

	.dataa(!Xd_0__inst_mult_10_488 ),
	.datab(!Xd_0__inst_mult_10_492 ),
	.datac(!Xd_0__inst_mult_10_496 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_337 ),
	.sharein(Xd_0__inst_mult_10_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_344 ),
	.cout(Xd_0__inst_mult_10_345 ),
	.shareout(Xd_0__inst_mult_10_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_111 (
// Equation(s):
// Xd_0__inst_mult_11_344  = SUM(( !Xd_0__inst_mult_11_484  $ (!Xd_0__inst_mult_11_488 ) ) + ( Xd_0__inst_mult_11_338  ) + ( Xd_0__inst_mult_11_337  ))
// Xd_0__inst_mult_11_345  = CARRY(( !Xd_0__inst_mult_11_484  $ (!Xd_0__inst_mult_11_488 ) ) + ( Xd_0__inst_mult_11_338  ) + ( Xd_0__inst_mult_11_337  ))
// Xd_0__inst_mult_11_346  = SHARE((Xd_0__inst_mult_11_484  & Xd_0__inst_mult_11_488 ))

	.dataa(!Xd_0__inst_mult_11_484 ),
	.datab(!Xd_0__inst_mult_11_488 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_337 ),
	.sharein(Xd_0__inst_mult_11_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_344 ),
	.cout(Xd_0__inst_mult_11_345 ),
	.shareout(Xd_0__inst_mult_11_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_112 (
// Equation(s):
// Xd_0__inst_mult_11_348  = SUM(( !Xd_0__inst_mult_11_492  $ (!Xd_0__inst_mult_11_496  $ (Xd_0__inst_mult_11_500 )) ) + ( Xd_0__inst_mult_11_342  ) + ( Xd_0__inst_mult_11_341  ))
// Xd_0__inst_mult_11_349  = CARRY(( !Xd_0__inst_mult_11_492  $ (!Xd_0__inst_mult_11_496  $ (Xd_0__inst_mult_11_500 )) ) + ( Xd_0__inst_mult_11_342  ) + ( Xd_0__inst_mult_11_341  ))
// Xd_0__inst_mult_11_350  = SHARE((!Xd_0__inst_mult_11_492  & (Xd_0__inst_mult_11_496  & Xd_0__inst_mult_11_500 )) # (Xd_0__inst_mult_11_492  & ((Xd_0__inst_mult_11_500 ) # (Xd_0__inst_mult_11_496 ))))

	.dataa(!Xd_0__inst_mult_11_492 ),
	.datab(!Xd_0__inst_mult_11_496 ),
	.datac(!Xd_0__inst_mult_11_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_341 ),
	.sharein(Xd_0__inst_mult_11_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_348 ),
	.cout(Xd_0__inst_mult_11_349 ),
	.shareout(Xd_0__inst_mult_11_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_111 (
// Equation(s):
// Xd_0__inst_mult_8_344  = SUM(( !Xd_0__inst_mult_8_484  $ (!Xd_0__inst_mult_8_488 ) ) + ( Xd_0__inst_mult_8_338  ) + ( Xd_0__inst_mult_8_337  ))
// Xd_0__inst_mult_8_345  = CARRY(( !Xd_0__inst_mult_8_484  $ (!Xd_0__inst_mult_8_488 ) ) + ( Xd_0__inst_mult_8_338  ) + ( Xd_0__inst_mult_8_337  ))
// Xd_0__inst_mult_8_346  = SHARE((Xd_0__inst_mult_8_484  & Xd_0__inst_mult_8_488 ))

	.dataa(!Xd_0__inst_mult_8_484 ),
	.datab(!Xd_0__inst_mult_8_488 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_337 ),
	.sharein(Xd_0__inst_mult_8_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_344 ),
	.cout(Xd_0__inst_mult_8_345 ),
	.shareout(Xd_0__inst_mult_8_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_112 (
// Equation(s):
// Xd_0__inst_mult_8_348  = SUM(( !Xd_0__inst_mult_8_492  $ (!Xd_0__inst_mult_8_496  $ (Xd_0__inst_mult_8_500 )) ) + ( Xd_0__inst_mult_8_342  ) + ( Xd_0__inst_mult_8_341  ))
// Xd_0__inst_mult_8_349  = CARRY(( !Xd_0__inst_mult_8_492  $ (!Xd_0__inst_mult_8_496  $ (Xd_0__inst_mult_8_500 )) ) + ( Xd_0__inst_mult_8_342  ) + ( Xd_0__inst_mult_8_341  ))
// Xd_0__inst_mult_8_350  = SHARE((!Xd_0__inst_mult_8_492  & (Xd_0__inst_mult_8_496  & Xd_0__inst_mult_8_500 )) # (Xd_0__inst_mult_8_492  & ((Xd_0__inst_mult_8_500 ) # (Xd_0__inst_mult_8_496 ))))

	.dataa(!Xd_0__inst_mult_8_492 ),
	.datab(!Xd_0__inst_mult_8_496 ),
	.datac(!Xd_0__inst_mult_8_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_341 ),
	.sharein(Xd_0__inst_mult_8_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_348 ),
	.cout(Xd_0__inst_mult_8_349 ),
	.shareout(Xd_0__inst_mult_8_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_107 (
// Equation(s):
// Xd_0__inst_mult_9_340  = SUM(( !Xd_0__inst_mult_9_480  $ (!Xd_0__inst_mult_9_484 ) ) + ( Xd_0__inst_mult_9_334  ) + ( Xd_0__inst_mult_9_333  ))
// Xd_0__inst_mult_9_341  = CARRY(( !Xd_0__inst_mult_9_480  $ (!Xd_0__inst_mult_9_484 ) ) + ( Xd_0__inst_mult_9_334  ) + ( Xd_0__inst_mult_9_333  ))
// Xd_0__inst_mult_9_342  = SHARE((Xd_0__inst_mult_9_480  & Xd_0__inst_mult_9_484 ))

	.dataa(!Xd_0__inst_mult_9_480 ),
	.datab(!Xd_0__inst_mult_9_484 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_333 ),
	.sharein(Xd_0__inst_mult_9_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_340 ),
	.cout(Xd_0__inst_mult_9_341 ),
	.shareout(Xd_0__inst_mult_9_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_108 (
// Equation(s):
// Xd_0__inst_mult_9_344  = SUM(( !Xd_0__inst_mult_9_488  $ (!Xd_0__inst_mult_9_492  $ (Xd_0__inst_mult_9_496 )) ) + ( Xd_0__inst_mult_9_338  ) + ( Xd_0__inst_mult_9_337  ))
// Xd_0__inst_mult_9_345  = CARRY(( !Xd_0__inst_mult_9_488  $ (!Xd_0__inst_mult_9_492  $ (Xd_0__inst_mult_9_496 )) ) + ( Xd_0__inst_mult_9_338  ) + ( Xd_0__inst_mult_9_337  ))
// Xd_0__inst_mult_9_346  = SHARE((!Xd_0__inst_mult_9_488  & (Xd_0__inst_mult_9_492  & Xd_0__inst_mult_9_496 )) # (Xd_0__inst_mult_9_488  & ((Xd_0__inst_mult_9_496 ) # (Xd_0__inst_mult_9_492 ))))

	.dataa(!Xd_0__inst_mult_9_488 ),
	.datab(!Xd_0__inst_mult_9_492 ),
	.datac(!Xd_0__inst_mult_9_496 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_337 ),
	.sharein(Xd_0__inst_mult_9_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_344 ),
	.cout(Xd_0__inst_mult_9_345 ),
	.shareout(Xd_0__inst_mult_9_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_107 (
// Equation(s):
// Xd_0__inst_mult_6_340  = SUM(( !Xd_0__inst_mult_6_480  $ (!Xd_0__inst_mult_6_484 ) ) + ( Xd_0__inst_mult_6_334  ) + ( Xd_0__inst_mult_6_333  ))
// Xd_0__inst_mult_6_341  = CARRY(( !Xd_0__inst_mult_6_480  $ (!Xd_0__inst_mult_6_484 ) ) + ( Xd_0__inst_mult_6_334  ) + ( Xd_0__inst_mult_6_333  ))
// Xd_0__inst_mult_6_342  = SHARE((Xd_0__inst_mult_6_480  & Xd_0__inst_mult_6_484 ))

	.dataa(!Xd_0__inst_mult_6_480 ),
	.datab(!Xd_0__inst_mult_6_484 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_333 ),
	.sharein(Xd_0__inst_mult_6_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_340 ),
	.cout(Xd_0__inst_mult_6_341 ),
	.shareout(Xd_0__inst_mult_6_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_108 (
// Equation(s):
// Xd_0__inst_mult_6_344  = SUM(( !Xd_0__inst_mult_6_488  $ (!Xd_0__inst_mult_6_492  $ (Xd_0__inst_mult_6_496 )) ) + ( Xd_0__inst_mult_6_338  ) + ( Xd_0__inst_mult_6_337  ))
// Xd_0__inst_mult_6_345  = CARRY(( !Xd_0__inst_mult_6_488  $ (!Xd_0__inst_mult_6_492  $ (Xd_0__inst_mult_6_496 )) ) + ( Xd_0__inst_mult_6_338  ) + ( Xd_0__inst_mult_6_337  ))
// Xd_0__inst_mult_6_346  = SHARE((!Xd_0__inst_mult_6_488  & (Xd_0__inst_mult_6_492  & Xd_0__inst_mult_6_496 )) # (Xd_0__inst_mult_6_488  & ((Xd_0__inst_mult_6_496 ) # (Xd_0__inst_mult_6_492 ))))

	.dataa(!Xd_0__inst_mult_6_488 ),
	.datab(!Xd_0__inst_mult_6_492 ),
	.datac(!Xd_0__inst_mult_6_496 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_337 ),
	.sharein(Xd_0__inst_mult_6_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_344 ),
	.cout(Xd_0__inst_mult_6_345 ),
	.shareout(Xd_0__inst_mult_6_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_101 (
// Equation(s):
// Xd_0__inst_mult_7_316  = SUM(( !Xd_0__inst_mult_7_464  $ (!Xd_0__inst_mult_7_468 ) ) + ( Xd_0__inst_mult_7_310  ) + ( Xd_0__inst_mult_7_309  ))
// Xd_0__inst_mult_7_317  = CARRY(( !Xd_0__inst_mult_7_464  $ (!Xd_0__inst_mult_7_468 ) ) + ( Xd_0__inst_mult_7_310  ) + ( Xd_0__inst_mult_7_309  ))
// Xd_0__inst_mult_7_318  = SHARE((Xd_0__inst_mult_7_464  & Xd_0__inst_mult_7_468 ))

	.dataa(!Xd_0__inst_mult_7_464 ),
	.datab(!Xd_0__inst_mult_7_468 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_309 ),
	.sharein(Xd_0__inst_mult_7_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_316 ),
	.cout(Xd_0__inst_mult_7_317 ),
	.shareout(Xd_0__inst_mult_7_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_102 (
// Equation(s):
// Xd_0__inst_mult_7_320  = SUM(( !Xd_0__inst_mult_7_472  $ (!Xd_0__inst_mult_7_476  $ (Xd_0__inst_mult_7_480 )) ) + ( Xd_0__inst_mult_7_314  ) + ( Xd_0__inst_mult_7_313  ))
// Xd_0__inst_mult_7_321  = CARRY(( !Xd_0__inst_mult_7_472  $ (!Xd_0__inst_mult_7_476  $ (Xd_0__inst_mult_7_480 )) ) + ( Xd_0__inst_mult_7_314  ) + ( Xd_0__inst_mult_7_313  ))
// Xd_0__inst_mult_7_322  = SHARE((!Xd_0__inst_mult_7_472  & (Xd_0__inst_mult_7_476  & Xd_0__inst_mult_7_480 )) # (Xd_0__inst_mult_7_472  & ((Xd_0__inst_mult_7_480 ) # (Xd_0__inst_mult_7_476 ))))

	.dataa(!Xd_0__inst_mult_7_472 ),
	.datab(!Xd_0__inst_mult_7_476 ),
	.datac(!Xd_0__inst_mult_7_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_313 ),
	.sharein(Xd_0__inst_mult_7_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_320 ),
	.cout(Xd_0__inst_mult_7_321 ),
	.shareout(Xd_0__inst_mult_7_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_113 (
// Equation(s):
// Xd_0__inst_mult_4_352  = SUM(( !Xd_0__inst_mult_4_504  $ (!Xd_0__inst_mult_4_508 ) ) + ( Xd_0__inst_mult_4_346  ) + ( Xd_0__inst_mult_4_345  ))
// Xd_0__inst_mult_4_353  = CARRY(( !Xd_0__inst_mult_4_504  $ (!Xd_0__inst_mult_4_508 ) ) + ( Xd_0__inst_mult_4_346  ) + ( Xd_0__inst_mult_4_345  ))
// Xd_0__inst_mult_4_354  = SHARE((Xd_0__inst_mult_4_504  & Xd_0__inst_mult_4_508 ))

	.dataa(!Xd_0__inst_mult_4_504 ),
	.datab(!Xd_0__inst_mult_4_508 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_345 ),
	.sharein(Xd_0__inst_mult_4_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_352 ),
	.cout(Xd_0__inst_mult_4_353 ),
	.shareout(Xd_0__inst_mult_4_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_114 (
// Equation(s):
// Xd_0__inst_mult_4_356  = SUM(( !Xd_0__inst_mult_4_512  $ (!Xd_0__inst_mult_4_412  $ (Xd_0__inst_mult_4_516 )) ) + ( Xd_0__inst_mult_4_350  ) + ( Xd_0__inst_mult_4_349  ))
// Xd_0__inst_mult_4_357  = CARRY(( !Xd_0__inst_mult_4_512  $ (!Xd_0__inst_mult_4_412  $ (Xd_0__inst_mult_4_516 )) ) + ( Xd_0__inst_mult_4_350  ) + ( Xd_0__inst_mult_4_349  ))
// Xd_0__inst_mult_4_358  = SHARE((!Xd_0__inst_mult_4_512  & (Xd_0__inst_mult_4_412  & Xd_0__inst_mult_4_516 )) # (Xd_0__inst_mult_4_512  & ((Xd_0__inst_mult_4_516 ) # (Xd_0__inst_mult_4_412 ))))

	.dataa(!Xd_0__inst_mult_4_512 ),
	.datab(!Xd_0__inst_mult_4_412 ),
	.datac(!Xd_0__inst_mult_4_516 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_349 ),
	.sharein(Xd_0__inst_mult_4_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_356 ),
	.cout(Xd_0__inst_mult_4_357 ),
	.shareout(Xd_0__inst_mult_4_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_101 (
// Equation(s):
// Xd_0__inst_mult_5_316  = SUM(( !Xd_0__inst_mult_5_464  $ (!Xd_0__inst_mult_5_468 ) ) + ( Xd_0__inst_mult_5_310  ) + ( Xd_0__inst_mult_5_309  ))
// Xd_0__inst_mult_5_317  = CARRY(( !Xd_0__inst_mult_5_464  $ (!Xd_0__inst_mult_5_468 ) ) + ( Xd_0__inst_mult_5_310  ) + ( Xd_0__inst_mult_5_309  ))
// Xd_0__inst_mult_5_318  = SHARE((Xd_0__inst_mult_5_464  & Xd_0__inst_mult_5_468 ))

	.dataa(!Xd_0__inst_mult_5_464 ),
	.datab(!Xd_0__inst_mult_5_468 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_309 ),
	.sharein(Xd_0__inst_mult_5_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_316 ),
	.cout(Xd_0__inst_mult_5_317 ),
	.shareout(Xd_0__inst_mult_5_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_102 (
// Equation(s):
// Xd_0__inst_mult_5_320  = SUM(( !Xd_0__inst_mult_5_472  $ (!Xd_0__inst_mult_5_476  $ (Xd_0__inst_mult_5_480 )) ) + ( Xd_0__inst_mult_5_314  ) + ( Xd_0__inst_mult_5_313  ))
// Xd_0__inst_mult_5_321  = CARRY(( !Xd_0__inst_mult_5_472  $ (!Xd_0__inst_mult_5_476  $ (Xd_0__inst_mult_5_480 )) ) + ( Xd_0__inst_mult_5_314  ) + ( Xd_0__inst_mult_5_313  ))
// Xd_0__inst_mult_5_322  = SHARE((!Xd_0__inst_mult_5_472  & (Xd_0__inst_mult_5_476  & Xd_0__inst_mult_5_480 )) # (Xd_0__inst_mult_5_472  & ((Xd_0__inst_mult_5_480 ) # (Xd_0__inst_mult_5_476 ))))

	.dataa(!Xd_0__inst_mult_5_472 ),
	.datab(!Xd_0__inst_mult_5_476 ),
	.datac(!Xd_0__inst_mult_5_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_313 ),
	.sharein(Xd_0__inst_mult_5_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_320 ),
	.cout(Xd_0__inst_mult_5_321 ),
	.shareout(Xd_0__inst_mult_5_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_105 (
// Equation(s):
// Xd_0__inst_mult_2_320  = SUM(( !Xd_0__inst_mult_2_468  $ (!Xd_0__inst_mult_2_472 ) ) + ( Xd_0__inst_mult_2_314  ) + ( Xd_0__inst_mult_2_313  ))
// Xd_0__inst_mult_2_321  = CARRY(( !Xd_0__inst_mult_2_468  $ (!Xd_0__inst_mult_2_472 ) ) + ( Xd_0__inst_mult_2_314  ) + ( Xd_0__inst_mult_2_313  ))
// Xd_0__inst_mult_2_322  = SHARE((Xd_0__inst_mult_2_468  & Xd_0__inst_mult_2_472 ))

	.dataa(!Xd_0__inst_mult_2_468 ),
	.datab(!Xd_0__inst_mult_2_472 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_313 ),
	.sharein(Xd_0__inst_mult_2_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_320 ),
	.cout(Xd_0__inst_mult_2_321 ),
	.shareout(Xd_0__inst_mult_2_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_106 (
// Equation(s):
// Xd_0__inst_mult_2_324  = SUM(( !Xd_0__inst_mult_2_476  $ (!Xd_0__inst_mult_2_480  $ (Xd_0__inst_mult_2_484 )) ) + ( Xd_0__inst_mult_2_318  ) + ( Xd_0__inst_mult_2_317  ))
// Xd_0__inst_mult_2_325  = CARRY(( !Xd_0__inst_mult_2_476  $ (!Xd_0__inst_mult_2_480  $ (Xd_0__inst_mult_2_484 )) ) + ( Xd_0__inst_mult_2_318  ) + ( Xd_0__inst_mult_2_317  ))
// Xd_0__inst_mult_2_326  = SHARE((!Xd_0__inst_mult_2_476  & (Xd_0__inst_mult_2_480  & Xd_0__inst_mult_2_484 )) # (Xd_0__inst_mult_2_476  & ((Xd_0__inst_mult_2_484 ) # (Xd_0__inst_mult_2_480 ))))

	.dataa(!Xd_0__inst_mult_2_476 ),
	.datab(!Xd_0__inst_mult_2_480 ),
	.datac(!Xd_0__inst_mult_2_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_317 ),
	.sharein(Xd_0__inst_mult_2_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_324 ),
	.cout(Xd_0__inst_mult_2_325 ),
	.shareout(Xd_0__inst_mult_2_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_101 (
// Equation(s):
// Xd_0__inst_mult_3_316  = SUM(( !Xd_0__inst_mult_3_464  $ (!Xd_0__inst_mult_3_468 ) ) + ( Xd_0__inst_mult_3_310  ) + ( Xd_0__inst_mult_3_309  ))
// Xd_0__inst_mult_3_317  = CARRY(( !Xd_0__inst_mult_3_464  $ (!Xd_0__inst_mult_3_468 ) ) + ( Xd_0__inst_mult_3_310  ) + ( Xd_0__inst_mult_3_309  ))
// Xd_0__inst_mult_3_318  = SHARE((Xd_0__inst_mult_3_464  & Xd_0__inst_mult_3_468 ))

	.dataa(!Xd_0__inst_mult_3_464 ),
	.datab(!Xd_0__inst_mult_3_468 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_309 ),
	.sharein(Xd_0__inst_mult_3_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_316 ),
	.cout(Xd_0__inst_mult_3_317 ),
	.shareout(Xd_0__inst_mult_3_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_102 (
// Equation(s):
// Xd_0__inst_mult_3_320  = SUM(( !Xd_0__inst_mult_3_472  $ (!Xd_0__inst_mult_3_476  $ (Xd_0__inst_mult_3_480 )) ) + ( Xd_0__inst_mult_3_314  ) + ( Xd_0__inst_mult_3_313  ))
// Xd_0__inst_mult_3_321  = CARRY(( !Xd_0__inst_mult_3_472  $ (!Xd_0__inst_mult_3_476  $ (Xd_0__inst_mult_3_480 )) ) + ( Xd_0__inst_mult_3_314  ) + ( Xd_0__inst_mult_3_313  ))
// Xd_0__inst_mult_3_322  = SHARE((!Xd_0__inst_mult_3_472  & (Xd_0__inst_mult_3_476  & Xd_0__inst_mult_3_480 )) # (Xd_0__inst_mult_3_472  & ((Xd_0__inst_mult_3_480 ) # (Xd_0__inst_mult_3_476 ))))

	.dataa(!Xd_0__inst_mult_3_472 ),
	.datab(!Xd_0__inst_mult_3_476 ),
	.datac(!Xd_0__inst_mult_3_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_313 ),
	.sharein(Xd_0__inst_mult_3_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_320 ),
	.cout(Xd_0__inst_mult_3_321 ),
	.shareout(Xd_0__inst_mult_3_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_105 (
// Equation(s):
// Xd_0__inst_mult_0_320  = SUM(( !Xd_0__inst_mult_0_468  $ (!Xd_0__inst_mult_0_472 ) ) + ( Xd_0__inst_mult_0_314  ) + ( Xd_0__inst_mult_0_313  ))
// Xd_0__inst_mult_0_321  = CARRY(( !Xd_0__inst_mult_0_468  $ (!Xd_0__inst_mult_0_472 ) ) + ( Xd_0__inst_mult_0_314  ) + ( Xd_0__inst_mult_0_313  ))
// Xd_0__inst_mult_0_322  = SHARE((Xd_0__inst_mult_0_468  & Xd_0__inst_mult_0_472 ))

	.dataa(!Xd_0__inst_mult_0_468 ),
	.datab(!Xd_0__inst_mult_0_472 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_313 ),
	.sharein(Xd_0__inst_mult_0_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_320 ),
	.cout(Xd_0__inst_mult_0_321 ),
	.shareout(Xd_0__inst_mult_0_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_106 (
// Equation(s):
// Xd_0__inst_mult_0_324  = SUM(( !Xd_0__inst_mult_0_476  $ (!Xd_0__inst_mult_0_480  $ (Xd_0__inst_mult_0_484 )) ) + ( Xd_0__inst_mult_0_318  ) + ( Xd_0__inst_mult_0_317  ))
// Xd_0__inst_mult_0_325  = CARRY(( !Xd_0__inst_mult_0_476  $ (!Xd_0__inst_mult_0_480  $ (Xd_0__inst_mult_0_484 )) ) + ( Xd_0__inst_mult_0_318  ) + ( Xd_0__inst_mult_0_317  ))
// Xd_0__inst_mult_0_326  = SHARE((!Xd_0__inst_mult_0_476  & (Xd_0__inst_mult_0_480  & Xd_0__inst_mult_0_484 )) # (Xd_0__inst_mult_0_476  & ((Xd_0__inst_mult_0_484 ) # (Xd_0__inst_mult_0_480 ))))

	.dataa(!Xd_0__inst_mult_0_476 ),
	.datab(!Xd_0__inst_mult_0_480 ),
	.datac(!Xd_0__inst_mult_0_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_317 ),
	.sharein(Xd_0__inst_mult_0_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_324 ),
	.cout(Xd_0__inst_mult_0_325 ),
	.shareout(Xd_0__inst_mult_0_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_105 (
// Equation(s):
// Xd_0__inst_mult_1_320  = SUM(( !Xd_0__inst_mult_1_468  $ (!Xd_0__inst_mult_1_472 ) ) + ( Xd_0__inst_mult_1_314  ) + ( Xd_0__inst_mult_1_313  ))
// Xd_0__inst_mult_1_321  = CARRY(( !Xd_0__inst_mult_1_468  $ (!Xd_0__inst_mult_1_472 ) ) + ( Xd_0__inst_mult_1_314  ) + ( Xd_0__inst_mult_1_313  ))
// Xd_0__inst_mult_1_322  = SHARE((Xd_0__inst_mult_1_468  & Xd_0__inst_mult_1_472 ))

	.dataa(!Xd_0__inst_mult_1_468 ),
	.datab(!Xd_0__inst_mult_1_472 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_313 ),
	.sharein(Xd_0__inst_mult_1_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_320 ),
	.cout(Xd_0__inst_mult_1_321 ),
	.shareout(Xd_0__inst_mult_1_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_106 (
// Equation(s):
// Xd_0__inst_mult_1_324  = SUM(( !Xd_0__inst_mult_1_476  $ (!Xd_0__inst_mult_1_480  $ (Xd_0__inst_mult_1_484 )) ) + ( Xd_0__inst_mult_1_318  ) + ( Xd_0__inst_mult_1_317  ))
// Xd_0__inst_mult_1_325  = CARRY(( !Xd_0__inst_mult_1_476  $ (!Xd_0__inst_mult_1_480  $ (Xd_0__inst_mult_1_484 )) ) + ( Xd_0__inst_mult_1_318  ) + ( Xd_0__inst_mult_1_317  ))
// Xd_0__inst_mult_1_326  = SHARE((!Xd_0__inst_mult_1_476  & (Xd_0__inst_mult_1_480  & Xd_0__inst_mult_1_484 )) # (Xd_0__inst_mult_1_476  & ((Xd_0__inst_mult_1_484 ) # (Xd_0__inst_mult_1_480 ))))

	.dataa(!Xd_0__inst_mult_1_476 ),
	.datab(!Xd_0__inst_mult_1_480 ),
	.datac(!Xd_0__inst_mult_1_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_317 ),
	.sharein(Xd_0__inst_mult_1_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_324 ),
	.cout(Xd_0__inst_mult_1_325 ),
	.shareout(Xd_0__inst_mult_1_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_115 (
// Equation(s):
// Xd_0__inst_mult_12_372  = SUM(( !Xd_0__inst_mult_12_528  $ (!Xd_0__inst_mult_12_532  $ (Xd_0__inst_mult_12_536 )) ) + ( Xd_0__inst_mult_12_370  ) + ( Xd_0__inst_mult_12_369  ))
// Xd_0__inst_mult_12_373  = CARRY(( !Xd_0__inst_mult_12_528  $ (!Xd_0__inst_mult_12_532  $ (Xd_0__inst_mult_12_536 )) ) + ( Xd_0__inst_mult_12_370  ) + ( Xd_0__inst_mult_12_369  ))
// Xd_0__inst_mult_12_374  = SHARE((!Xd_0__inst_mult_12_528  & (Xd_0__inst_mult_12_532  & Xd_0__inst_mult_12_536 )) # (Xd_0__inst_mult_12_528  & ((Xd_0__inst_mult_12_536 ) # (Xd_0__inst_mult_12_532 ))))

	.dataa(!Xd_0__inst_mult_12_528 ),
	.datab(!Xd_0__inst_mult_12_532 ),
	.datac(!Xd_0__inst_mult_12_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_369 ),
	.sharein(Xd_0__inst_mult_12_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_372 ),
	.cout(Xd_0__inst_mult_12_373 ),
	.shareout(Xd_0__inst_mult_12_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_113 (
// Equation(s):
// Xd_0__inst_mult_13_352  = SUM(( !Xd_0__inst_mult_13_504  $ (!Xd_0__inst_mult_13_508  $ (Xd_0__inst_mult_13_512 )) ) + ( Xd_0__inst_mult_13_350  ) + ( Xd_0__inst_mult_13_349  ))
// Xd_0__inst_mult_13_353  = CARRY(( !Xd_0__inst_mult_13_504  $ (!Xd_0__inst_mult_13_508  $ (Xd_0__inst_mult_13_512 )) ) + ( Xd_0__inst_mult_13_350  ) + ( Xd_0__inst_mult_13_349  ))
// Xd_0__inst_mult_13_354  = SHARE((!Xd_0__inst_mult_13_504  & (Xd_0__inst_mult_13_508  & Xd_0__inst_mult_13_512 )) # (Xd_0__inst_mult_13_504  & ((Xd_0__inst_mult_13_512 ) # (Xd_0__inst_mult_13_508 ))))

	.dataa(!Xd_0__inst_mult_13_504 ),
	.datab(!Xd_0__inst_mult_13_508 ),
	.datac(!Xd_0__inst_mult_13_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_349 ),
	.sharein(Xd_0__inst_mult_13_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_352 ),
	.cout(Xd_0__inst_mult_13_353 ),
	.shareout(Xd_0__inst_mult_13_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_117 (
// Equation(s):
// Xd_0__inst_mult_14_368  = SUM(( !Xd_0__inst_mult_14_504  $ (!Xd_0__inst_mult_14_508  $ (Xd_0__inst_mult_14_512 )) ) + ( Xd_0__inst_mult_14_366  ) + ( Xd_0__inst_mult_14_365  ))
// Xd_0__inst_mult_14_369  = CARRY(( !Xd_0__inst_mult_14_504  $ (!Xd_0__inst_mult_14_508  $ (Xd_0__inst_mult_14_512 )) ) + ( Xd_0__inst_mult_14_366  ) + ( Xd_0__inst_mult_14_365  ))
// Xd_0__inst_mult_14_370  = SHARE((!Xd_0__inst_mult_14_504  & (Xd_0__inst_mult_14_508  & Xd_0__inst_mult_14_512 )) # (Xd_0__inst_mult_14_504  & ((Xd_0__inst_mult_14_512 ) # (Xd_0__inst_mult_14_508 ))))

	.dataa(!Xd_0__inst_mult_14_504 ),
	.datab(!Xd_0__inst_mult_14_508 ),
	.datac(!Xd_0__inst_mult_14_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_365 ),
	.sharein(Xd_0__inst_mult_14_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_368 ),
	.cout(Xd_0__inst_mult_14_369 ),
	.shareout(Xd_0__inst_mult_14_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_119 (
// Equation(s):
// Xd_0__inst_mult_15_376  = SUM(( !Xd_0__inst_mult_15_532  $ (!Xd_0__inst_mult_15_536  $ (Xd_0__inst_mult_15_540 )) ) + ( Xd_0__inst_mult_15_374  ) + ( Xd_0__inst_mult_15_373  ))
// Xd_0__inst_mult_15_377  = CARRY(( !Xd_0__inst_mult_15_532  $ (!Xd_0__inst_mult_15_536  $ (Xd_0__inst_mult_15_540 )) ) + ( Xd_0__inst_mult_15_374  ) + ( Xd_0__inst_mult_15_373  ))
// Xd_0__inst_mult_15_378  = SHARE((!Xd_0__inst_mult_15_532  & (Xd_0__inst_mult_15_536  & Xd_0__inst_mult_15_540 )) # (Xd_0__inst_mult_15_532  & ((Xd_0__inst_mult_15_540 ) # (Xd_0__inst_mult_15_536 ))))

	.dataa(!Xd_0__inst_mult_15_532 ),
	.datab(!Xd_0__inst_mult_15_536 ),
	.datac(!Xd_0__inst_mult_15_540 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_373 ),
	.sharein(Xd_0__inst_mult_15_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_376 ),
	.cout(Xd_0__inst_mult_15_377 ),
	.shareout(Xd_0__inst_mult_15_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_109 (
// Equation(s):
// Xd_0__inst_mult_10_348  = SUM(( !Xd_0__inst_mult_10_500  $ (!Xd_0__inst_mult_10_504  $ (Xd_0__inst_mult_10_508 )) ) + ( Xd_0__inst_mult_10_346  ) + ( Xd_0__inst_mult_10_345  ))
// Xd_0__inst_mult_10_349  = CARRY(( !Xd_0__inst_mult_10_500  $ (!Xd_0__inst_mult_10_504  $ (Xd_0__inst_mult_10_508 )) ) + ( Xd_0__inst_mult_10_346  ) + ( Xd_0__inst_mult_10_345  ))
// Xd_0__inst_mult_10_350  = SHARE((!Xd_0__inst_mult_10_500  & (Xd_0__inst_mult_10_504  & Xd_0__inst_mult_10_508 )) # (Xd_0__inst_mult_10_500  & ((Xd_0__inst_mult_10_508 ) # (Xd_0__inst_mult_10_504 ))))

	.dataa(!Xd_0__inst_mult_10_500 ),
	.datab(!Xd_0__inst_mult_10_504 ),
	.datac(!Xd_0__inst_mult_10_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_345 ),
	.sharein(Xd_0__inst_mult_10_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_348 ),
	.cout(Xd_0__inst_mult_10_349 ),
	.shareout(Xd_0__inst_mult_10_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_113 (
// Equation(s):
// Xd_0__inst_mult_11_352  = SUM(( !Xd_0__inst_mult_11_504  $ (!Xd_0__inst_mult_11_508  $ (Xd_0__inst_mult_11_512 )) ) + ( Xd_0__inst_mult_11_350  ) + ( Xd_0__inst_mult_11_349  ))
// Xd_0__inst_mult_11_353  = CARRY(( !Xd_0__inst_mult_11_504  $ (!Xd_0__inst_mult_11_508  $ (Xd_0__inst_mult_11_512 )) ) + ( Xd_0__inst_mult_11_350  ) + ( Xd_0__inst_mult_11_349  ))
// Xd_0__inst_mult_11_354  = SHARE((!Xd_0__inst_mult_11_504  & (Xd_0__inst_mult_11_508  & Xd_0__inst_mult_11_512 )) # (Xd_0__inst_mult_11_504  & ((Xd_0__inst_mult_11_512 ) # (Xd_0__inst_mult_11_508 ))))

	.dataa(!Xd_0__inst_mult_11_504 ),
	.datab(!Xd_0__inst_mult_11_508 ),
	.datac(!Xd_0__inst_mult_11_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_349 ),
	.sharein(Xd_0__inst_mult_11_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_352 ),
	.cout(Xd_0__inst_mult_11_353 ),
	.shareout(Xd_0__inst_mult_11_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_113 (
// Equation(s):
// Xd_0__inst_mult_8_352  = SUM(( !Xd_0__inst_mult_8_504  $ (!Xd_0__inst_mult_8_508  $ (Xd_0__inst_mult_8_512 )) ) + ( Xd_0__inst_mult_8_350  ) + ( Xd_0__inst_mult_8_349  ))
// Xd_0__inst_mult_8_353  = CARRY(( !Xd_0__inst_mult_8_504  $ (!Xd_0__inst_mult_8_508  $ (Xd_0__inst_mult_8_512 )) ) + ( Xd_0__inst_mult_8_350  ) + ( Xd_0__inst_mult_8_349  ))
// Xd_0__inst_mult_8_354  = SHARE((!Xd_0__inst_mult_8_504  & (Xd_0__inst_mult_8_508  & Xd_0__inst_mult_8_512 )) # (Xd_0__inst_mult_8_504  & ((Xd_0__inst_mult_8_512 ) # (Xd_0__inst_mult_8_508 ))))

	.dataa(!Xd_0__inst_mult_8_504 ),
	.datab(!Xd_0__inst_mult_8_508 ),
	.datac(!Xd_0__inst_mult_8_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_349 ),
	.sharein(Xd_0__inst_mult_8_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_352 ),
	.cout(Xd_0__inst_mult_8_353 ),
	.shareout(Xd_0__inst_mult_8_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_109 (
// Equation(s):
// Xd_0__inst_mult_9_348  = SUM(( !Xd_0__inst_mult_9_500  $ (!Xd_0__inst_mult_9_504  $ (Xd_0__inst_mult_9_508 )) ) + ( Xd_0__inst_mult_9_346  ) + ( Xd_0__inst_mult_9_345  ))
// Xd_0__inst_mult_9_349  = CARRY(( !Xd_0__inst_mult_9_500  $ (!Xd_0__inst_mult_9_504  $ (Xd_0__inst_mult_9_508 )) ) + ( Xd_0__inst_mult_9_346  ) + ( Xd_0__inst_mult_9_345  ))
// Xd_0__inst_mult_9_350  = SHARE((!Xd_0__inst_mult_9_500  & (Xd_0__inst_mult_9_504  & Xd_0__inst_mult_9_508 )) # (Xd_0__inst_mult_9_500  & ((Xd_0__inst_mult_9_508 ) # (Xd_0__inst_mult_9_504 ))))

	.dataa(!Xd_0__inst_mult_9_500 ),
	.datab(!Xd_0__inst_mult_9_504 ),
	.datac(!Xd_0__inst_mult_9_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_345 ),
	.sharein(Xd_0__inst_mult_9_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_348 ),
	.cout(Xd_0__inst_mult_9_349 ),
	.shareout(Xd_0__inst_mult_9_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_109 (
// Equation(s):
// Xd_0__inst_mult_6_348  = SUM(( !Xd_0__inst_mult_6_500  $ (!Xd_0__inst_mult_6_504  $ (Xd_0__inst_mult_6_508 )) ) + ( Xd_0__inst_mult_6_346  ) + ( Xd_0__inst_mult_6_345  ))
// Xd_0__inst_mult_6_349  = CARRY(( !Xd_0__inst_mult_6_500  $ (!Xd_0__inst_mult_6_504  $ (Xd_0__inst_mult_6_508 )) ) + ( Xd_0__inst_mult_6_346  ) + ( Xd_0__inst_mult_6_345  ))
// Xd_0__inst_mult_6_350  = SHARE((!Xd_0__inst_mult_6_500  & (Xd_0__inst_mult_6_504  & Xd_0__inst_mult_6_508 )) # (Xd_0__inst_mult_6_500  & ((Xd_0__inst_mult_6_508 ) # (Xd_0__inst_mult_6_504 ))))

	.dataa(!Xd_0__inst_mult_6_500 ),
	.datab(!Xd_0__inst_mult_6_504 ),
	.datac(!Xd_0__inst_mult_6_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_345 ),
	.sharein(Xd_0__inst_mult_6_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_348 ),
	.cout(Xd_0__inst_mult_6_349 ),
	.shareout(Xd_0__inst_mult_6_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_103 (
// Equation(s):
// Xd_0__inst_mult_7_324  = SUM(( !Xd_0__inst_mult_7_484  $ (!Xd_0__inst_mult_7_488  $ (((din_b[86] & din_a[94])))) ) + ( Xd_0__inst_mult_7_318  ) + ( Xd_0__inst_mult_7_317  ))
// Xd_0__inst_mult_7_325  = CARRY(( !Xd_0__inst_mult_7_484  $ (!Xd_0__inst_mult_7_488  $ (((din_b[86] & din_a[94])))) ) + ( Xd_0__inst_mult_7_318  ) + ( Xd_0__inst_mult_7_317  ))
// Xd_0__inst_mult_7_326  = SHARE((!Xd_0__inst_mult_7_484  & (Xd_0__inst_mult_7_488  & (din_b[86] & din_a[94]))) # (Xd_0__inst_mult_7_484  & (((din_b[86] & din_a[94])) # (Xd_0__inst_mult_7_488 ))))

	.dataa(!Xd_0__inst_mult_7_484 ),
	.datab(!Xd_0__inst_mult_7_488 ),
	.datac(!din_b[86]),
	.datad(!din_a[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_317 ),
	.sharein(Xd_0__inst_mult_7_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_324 ),
	.cout(Xd_0__inst_mult_7_325 ),
	.shareout(Xd_0__inst_mult_7_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_104 (
// Equation(s):
// Xd_0__inst_mult_7_328  = SUM(( !Xd_0__inst_mult_7_492  $ (!Xd_0__inst_mult_7_496  $ (Xd_0__inst_mult_7_500 )) ) + ( Xd_0__inst_mult_7_322  ) + ( Xd_0__inst_mult_7_321  ))
// Xd_0__inst_mult_7_329  = CARRY(( !Xd_0__inst_mult_7_492  $ (!Xd_0__inst_mult_7_496  $ (Xd_0__inst_mult_7_500 )) ) + ( Xd_0__inst_mult_7_322  ) + ( Xd_0__inst_mult_7_321  ))
// Xd_0__inst_mult_7_330  = SHARE((!Xd_0__inst_mult_7_492  & (Xd_0__inst_mult_7_496  & Xd_0__inst_mult_7_500 )) # (Xd_0__inst_mult_7_492  & ((Xd_0__inst_mult_7_500 ) # (Xd_0__inst_mult_7_496 ))))

	.dataa(!Xd_0__inst_mult_7_492 ),
	.datab(!Xd_0__inst_mult_7_496 ),
	.datac(!Xd_0__inst_mult_7_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_321 ),
	.sharein(Xd_0__inst_mult_7_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_328 ),
	.cout(Xd_0__inst_mult_7_329 ),
	.shareout(Xd_0__inst_mult_7_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_115 (
// Equation(s):
// Xd_0__inst_mult_4_360  = SUM(( !Xd_0__inst_mult_4_520  $ (!Xd_0__inst_mult_4_524  $ (((din_b[50] & din_a[58])))) ) + ( Xd_0__inst_mult_4_354  ) + ( Xd_0__inst_mult_4_353  ))
// Xd_0__inst_mult_4_361  = CARRY(( !Xd_0__inst_mult_4_520  $ (!Xd_0__inst_mult_4_524  $ (((din_b[50] & din_a[58])))) ) + ( Xd_0__inst_mult_4_354  ) + ( Xd_0__inst_mult_4_353  ))
// Xd_0__inst_mult_4_362  = SHARE((!Xd_0__inst_mult_4_520  & (Xd_0__inst_mult_4_524  & (din_b[50] & din_a[58]))) # (Xd_0__inst_mult_4_520  & (((din_b[50] & din_a[58])) # (Xd_0__inst_mult_4_524 ))))

	.dataa(!Xd_0__inst_mult_4_520 ),
	.datab(!Xd_0__inst_mult_4_524 ),
	.datac(!din_b[50]),
	.datad(!din_a[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_353 ),
	.sharein(Xd_0__inst_mult_4_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_360 ),
	.cout(Xd_0__inst_mult_4_361 ),
	.shareout(Xd_0__inst_mult_4_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_116 (
// Equation(s):
// Xd_0__inst_mult_4_364  = SUM(( !Xd_0__inst_mult_4_528  $ (!Xd_0__inst_mult_4_288  $ (Xd_0__inst_mult_4_532 )) ) + ( Xd_0__inst_mult_4_358  ) + ( Xd_0__inst_mult_4_357  ))
// Xd_0__inst_mult_4_365  = CARRY(( !Xd_0__inst_mult_4_528  $ (!Xd_0__inst_mult_4_288  $ (Xd_0__inst_mult_4_532 )) ) + ( Xd_0__inst_mult_4_358  ) + ( Xd_0__inst_mult_4_357  ))
// Xd_0__inst_mult_4_366  = SHARE((!Xd_0__inst_mult_4_528  & (Xd_0__inst_mult_4_288  & Xd_0__inst_mult_4_532 )) # (Xd_0__inst_mult_4_528  & ((Xd_0__inst_mult_4_532 ) # (Xd_0__inst_mult_4_288 ))))

	.dataa(!Xd_0__inst_mult_4_528 ),
	.datab(!Xd_0__inst_mult_4_288 ),
	.datac(!Xd_0__inst_mult_4_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_357 ),
	.sharein(Xd_0__inst_mult_4_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_364 ),
	.cout(Xd_0__inst_mult_4_365 ),
	.shareout(Xd_0__inst_mult_4_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_103 (
// Equation(s):
// Xd_0__inst_mult_5_324  = SUM(( !Xd_0__inst_mult_5_484  $ (!Xd_0__inst_mult_5_488  $ (((din_b[62] & din_a[70])))) ) + ( Xd_0__inst_mult_5_318  ) + ( Xd_0__inst_mult_5_317  ))
// Xd_0__inst_mult_5_325  = CARRY(( !Xd_0__inst_mult_5_484  $ (!Xd_0__inst_mult_5_488  $ (((din_b[62] & din_a[70])))) ) + ( Xd_0__inst_mult_5_318  ) + ( Xd_0__inst_mult_5_317  ))
// Xd_0__inst_mult_5_326  = SHARE((!Xd_0__inst_mult_5_484  & (Xd_0__inst_mult_5_488  & (din_b[62] & din_a[70]))) # (Xd_0__inst_mult_5_484  & (((din_b[62] & din_a[70])) # (Xd_0__inst_mult_5_488 ))))

	.dataa(!Xd_0__inst_mult_5_484 ),
	.datab(!Xd_0__inst_mult_5_488 ),
	.datac(!din_b[62]),
	.datad(!din_a[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_317 ),
	.sharein(Xd_0__inst_mult_5_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_324 ),
	.cout(Xd_0__inst_mult_5_325 ),
	.shareout(Xd_0__inst_mult_5_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_104 (
// Equation(s):
// Xd_0__inst_mult_5_328  = SUM(( !Xd_0__inst_mult_5_492  $ (!Xd_0__inst_mult_5_496  $ (Xd_0__inst_mult_5_500 )) ) + ( Xd_0__inst_mult_5_322  ) + ( Xd_0__inst_mult_5_321  ))
// Xd_0__inst_mult_5_329  = CARRY(( !Xd_0__inst_mult_5_492  $ (!Xd_0__inst_mult_5_496  $ (Xd_0__inst_mult_5_500 )) ) + ( Xd_0__inst_mult_5_322  ) + ( Xd_0__inst_mult_5_321  ))
// Xd_0__inst_mult_5_330  = SHARE((!Xd_0__inst_mult_5_492  & (Xd_0__inst_mult_5_496  & Xd_0__inst_mult_5_500 )) # (Xd_0__inst_mult_5_492  & ((Xd_0__inst_mult_5_500 ) # (Xd_0__inst_mult_5_496 ))))

	.dataa(!Xd_0__inst_mult_5_492 ),
	.datab(!Xd_0__inst_mult_5_496 ),
	.datac(!Xd_0__inst_mult_5_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_321 ),
	.sharein(Xd_0__inst_mult_5_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_328 ),
	.cout(Xd_0__inst_mult_5_329 ),
	.shareout(Xd_0__inst_mult_5_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_107 (
// Equation(s):
// Xd_0__inst_mult_2_328  = SUM(( !Xd_0__inst_mult_2_488  $ (!Xd_0__inst_mult_2_492  $ (((din_b[26] & din_a[34])))) ) + ( Xd_0__inst_mult_2_322  ) + ( Xd_0__inst_mult_2_321  ))
// Xd_0__inst_mult_2_329  = CARRY(( !Xd_0__inst_mult_2_488  $ (!Xd_0__inst_mult_2_492  $ (((din_b[26] & din_a[34])))) ) + ( Xd_0__inst_mult_2_322  ) + ( Xd_0__inst_mult_2_321  ))
// Xd_0__inst_mult_2_330  = SHARE((!Xd_0__inst_mult_2_488  & (Xd_0__inst_mult_2_492  & (din_b[26] & din_a[34]))) # (Xd_0__inst_mult_2_488  & (((din_b[26] & din_a[34])) # (Xd_0__inst_mult_2_492 ))))

	.dataa(!Xd_0__inst_mult_2_488 ),
	.datab(!Xd_0__inst_mult_2_492 ),
	.datac(!din_b[26]),
	.datad(!din_a[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_321 ),
	.sharein(Xd_0__inst_mult_2_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_328 ),
	.cout(Xd_0__inst_mult_2_329 ),
	.shareout(Xd_0__inst_mult_2_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_108 (
// Equation(s):
// Xd_0__inst_mult_2_332  = SUM(( !Xd_0__inst_mult_2_496  $ (!Xd_0__inst_mult_2_500  $ (Xd_0__inst_mult_2_504 )) ) + ( Xd_0__inst_mult_2_326  ) + ( Xd_0__inst_mult_2_325  ))
// Xd_0__inst_mult_2_333  = CARRY(( !Xd_0__inst_mult_2_496  $ (!Xd_0__inst_mult_2_500  $ (Xd_0__inst_mult_2_504 )) ) + ( Xd_0__inst_mult_2_326  ) + ( Xd_0__inst_mult_2_325  ))
// Xd_0__inst_mult_2_334  = SHARE((!Xd_0__inst_mult_2_496  & (Xd_0__inst_mult_2_500  & Xd_0__inst_mult_2_504 )) # (Xd_0__inst_mult_2_496  & ((Xd_0__inst_mult_2_504 ) # (Xd_0__inst_mult_2_500 ))))

	.dataa(!Xd_0__inst_mult_2_496 ),
	.datab(!Xd_0__inst_mult_2_500 ),
	.datac(!Xd_0__inst_mult_2_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_325 ),
	.sharein(Xd_0__inst_mult_2_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_332 ),
	.cout(Xd_0__inst_mult_2_333 ),
	.shareout(Xd_0__inst_mult_2_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_103 (
// Equation(s):
// Xd_0__inst_mult_3_324  = SUM(( !Xd_0__inst_mult_3_484  $ (!Xd_0__inst_mult_3_488  $ (((din_b[38] & din_a[46])))) ) + ( Xd_0__inst_mult_3_318  ) + ( Xd_0__inst_mult_3_317  ))
// Xd_0__inst_mult_3_325  = CARRY(( !Xd_0__inst_mult_3_484  $ (!Xd_0__inst_mult_3_488  $ (((din_b[38] & din_a[46])))) ) + ( Xd_0__inst_mult_3_318  ) + ( Xd_0__inst_mult_3_317  ))
// Xd_0__inst_mult_3_326  = SHARE((!Xd_0__inst_mult_3_484  & (Xd_0__inst_mult_3_488  & (din_b[38] & din_a[46]))) # (Xd_0__inst_mult_3_484  & (((din_b[38] & din_a[46])) # (Xd_0__inst_mult_3_488 ))))

	.dataa(!Xd_0__inst_mult_3_484 ),
	.datab(!Xd_0__inst_mult_3_488 ),
	.datac(!din_b[38]),
	.datad(!din_a[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_317 ),
	.sharein(Xd_0__inst_mult_3_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_324 ),
	.cout(Xd_0__inst_mult_3_325 ),
	.shareout(Xd_0__inst_mult_3_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_104 (
// Equation(s):
// Xd_0__inst_mult_3_328  = SUM(( !Xd_0__inst_mult_3_492  $ (!Xd_0__inst_mult_3_496  $ (Xd_0__inst_mult_3_500 )) ) + ( Xd_0__inst_mult_3_322  ) + ( Xd_0__inst_mult_3_321  ))
// Xd_0__inst_mult_3_329  = CARRY(( !Xd_0__inst_mult_3_492  $ (!Xd_0__inst_mult_3_496  $ (Xd_0__inst_mult_3_500 )) ) + ( Xd_0__inst_mult_3_322  ) + ( Xd_0__inst_mult_3_321  ))
// Xd_0__inst_mult_3_330  = SHARE((!Xd_0__inst_mult_3_492  & (Xd_0__inst_mult_3_496  & Xd_0__inst_mult_3_500 )) # (Xd_0__inst_mult_3_492  & ((Xd_0__inst_mult_3_500 ) # (Xd_0__inst_mult_3_496 ))))

	.dataa(!Xd_0__inst_mult_3_492 ),
	.datab(!Xd_0__inst_mult_3_496 ),
	.datac(!Xd_0__inst_mult_3_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_321 ),
	.sharein(Xd_0__inst_mult_3_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_328 ),
	.cout(Xd_0__inst_mult_3_329 ),
	.shareout(Xd_0__inst_mult_3_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_107 (
// Equation(s):
// Xd_0__inst_mult_0_328  = SUM(( !Xd_0__inst_mult_0_488  $ (!Xd_0__inst_mult_0_492  $ (((din_b[2] & din_a[10])))) ) + ( Xd_0__inst_mult_0_322  ) + ( Xd_0__inst_mult_0_321  ))
// Xd_0__inst_mult_0_329  = CARRY(( !Xd_0__inst_mult_0_488  $ (!Xd_0__inst_mult_0_492  $ (((din_b[2] & din_a[10])))) ) + ( Xd_0__inst_mult_0_322  ) + ( Xd_0__inst_mult_0_321  ))
// Xd_0__inst_mult_0_330  = SHARE((!Xd_0__inst_mult_0_488  & (Xd_0__inst_mult_0_492  & (din_b[2] & din_a[10]))) # (Xd_0__inst_mult_0_488  & (((din_b[2] & din_a[10])) # (Xd_0__inst_mult_0_492 ))))

	.dataa(!Xd_0__inst_mult_0_488 ),
	.datab(!Xd_0__inst_mult_0_492 ),
	.datac(!din_b[2]),
	.datad(!din_a[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_321 ),
	.sharein(Xd_0__inst_mult_0_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_328 ),
	.cout(Xd_0__inst_mult_0_329 ),
	.shareout(Xd_0__inst_mult_0_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_108 (
// Equation(s):
// Xd_0__inst_mult_0_332  = SUM(( !Xd_0__inst_mult_0_496  $ (!Xd_0__inst_mult_0_500  $ (Xd_0__inst_mult_0_504 )) ) + ( Xd_0__inst_mult_0_326  ) + ( Xd_0__inst_mult_0_325  ))
// Xd_0__inst_mult_0_333  = CARRY(( !Xd_0__inst_mult_0_496  $ (!Xd_0__inst_mult_0_500  $ (Xd_0__inst_mult_0_504 )) ) + ( Xd_0__inst_mult_0_326  ) + ( Xd_0__inst_mult_0_325  ))
// Xd_0__inst_mult_0_334  = SHARE((!Xd_0__inst_mult_0_496  & (Xd_0__inst_mult_0_500  & Xd_0__inst_mult_0_504 )) # (Xd_0__inst_mult_0_496  & ((Xd_0__inst_mult_0_504 ) # (Xd_0__inst_mult_0_500 ))))

	.dataa(!Xd_0__inst_mult_0_496 ),
	.datab(!Xd_0__inst_mult_0_500 ),
	.datac(!Xd_0__inst_mult_0_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_325 ),
	.sharein(Xd_0__inst_mult_0_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_332 ),
	.cout(Xd_0__inst_mult_0_333 ),
	.shareout(Xd_0__inst_mult_0_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_107 (
// Equation(s):
// Xd_0__inst_mult_1_328  = SUM(( !Xd_0__inst_mult_1_488  $ (!Xd_0__inst_mult_1_492  $ (((din_b[14] & din_a[22])))) ) + ( Xd_0__inst_mult_1_322  ) + ( Xd_0__inst_mult_1_321  ))
// Xd_0__inst_mult_1_329  = CARRY(( !Xd_0__inst_mult_1_488  $ (!Xd_0__inst_mult_1_492  $ (((din_b[14] & din_a[22])))) ) + ( Xd_0__inst_mult_1_322  ) + ( Xd_0__inst_mult_1_321  ))
// Xd_0__inst_mult_1_330  = SHARE((!Xd_0__inst_mult_1_488  & (Xd_0__inst_mult_1_492  & (din_b[14] & din_a[22]))) # (Xd_0__inst_mult_1_488  & (((din_b[14] & din_a[22])) # (Xd_0__inst_mult_1_492 ))))

	.dataa(!Xd_0__inst_mult_1_488 ),
	.datab(!Xd_0__inst_mult_1_492 ),
	.datac(!din_b[14]),
	.datad(!din_a[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_321 ),
	.sharein(Xd_0__inst_mult_1_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_328 ),
	.cout(Xd_0__inst_mult_1_329 ),
	.shareout(Xd_0__inst_mult_1_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_108 (
// Equation(s):
// Xd_0__inst_mult_1_332  = SUM(( !Xd_0__inst_mult_1_496  $ (!Xd_0__inst_mult_1_500  $ (Xd_0__inst_mult_1_504 )) ) + ( Xd_0__inst_mult_1_326  ) + ( Xd_0__inst_mult_1_325  ))
// Xd_0__inst_mult_1_333  = CARRY(( !Xd_0__inst_mult_1_496  $ (!Xd_0__inst_mult_1_500  $ (Xd_0__inst_mult_1_504 )) ) + ( Xd_0__inst_mult_1_326  ) + ( Xd_0__inst_mult_1_325  ))
// Xd_0__inst_mult_1_334  = SHARE((!Xd_0__inst_mult_1_496  & (Xd_0__inst_mult_1_500  & Xd_0__inst_mult_1_504 )) # (Xd_0__inst_mult_1_496  & ((Xd_0__inst_mult_1_504 ) # (Xd_0__inst_mult_1_500 ))))

	.dataa(!Xd_0__inst_mult_1_496 ),
	.datab(!Xd_0__inst_mult_1_500 ),
	.datac(!Xd_0__inst_mult_1_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_325 ),
	.sharein(Xd_0__inst_mult_1_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_332 ),
	.cout(Xd_0__inst_mult_1_333 ),
	.shareout(Xd_0__inst_mult_1_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_116 (
// Equation(s):
// Xd_0__inst_mult_12_376  = SUM(( !Xd_0__inst_mult_12_540  $ (!Xd_0__inst_mult_12_416  $ (Xd_0__inst_mult_12_544 )) ) + ( Xd_0__inst_mult_12_374  ) + ( Xd_0__inst_mult_12_373  ))
// Xd_0__inst_mult_12_377  = CARRY(( !Xd_0__inst_mult_12_540  $ (!Xd_0__inst_mult_12_416  $ (Xd_0__inst_mult_12_544 )) ) + ( Xd_0__inst_mult_12_374  ) + ( Xd_0__inst_mult_12_373  ))
// Xd_0__inst_mult_12_378  = SHARE((!Xd_0__inst_mult_12_540  & (Xd_0__inst_mult_12_416  & Xd_0__inst_mult_12_544 )) # (Xd_0__inst_mult_12_540  & ((Xd_0__inst_mult_12_544 ) # (Xd_0__inst_mult_12_416 ))))

	.dataa(!Xd_0__inst_mult_12_540 ),
	.datab(!Xd_0__inst_mult_12_416 ),
	.datac(!Xd_0__inst_mult_12_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_373 ),
	.sharein(Xd_0__inst_mult_12_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_376 ),
	.cout(Xd_0__inst_mult_12_377 ),
	.shareout(Xd_0__inst_mult_12_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_114 (
// Equation(s):
// Xd_0__inst_mult_13_356  = SUM(( !Xd_0__inst_mult_13_516  $ (!Xd_0__inst_mult_13_520  $ (Xd_0__inst_mult_13_524 )) ) + ( Xd_0__inst_mult_13_354  ) + ( Xd_0__inst_mult_13_353  ))
// Xd_0__inst_mult_13_357  = CARRY(( !Xd_0__inst_mult_13_516  $ (!Xd_0__inst_mult_13_520  $ (Xd_0__inst_mult_13_524 )) ) + ( Xd_0__inst_mult_13_354  ) + ( Xd_0__inst_mult_13_353  ))
// Xd_0__inst_mult_13_358  = SHARE((!Xd_0__inst_mult_13_516  & (Xd_0__inst_mult_13_520  & Xd_0__inst_mult_13_524 )) # (Xd_0__inst_mult_13_516  & ((Xd_0__inst_mult_13_524 ) # (Xd_0__inst_mult_13_520 ))))

	.dataa(!Xd_0__inst_mult_13_516 ),
	.datab(!Xd_0__inst_mult_13_520 ),
	.datac(!Xd_0__inst_mult_13_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_353 ),
	.sharein(Xd_0__inst_mult_13_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_356 ),
	.cout(Xd_0__inst_mult_13_357 ),
	.shareout(Xd_0__inst_mult_13_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_118 (
// Equation(s):
// Xd_0__inst_mult_14_372  = SUM(( !Xd_0__inst_mult_14_516  $ (!Xd_0__inst_mult_14_520  $ (Xd_0__inst_mult_14_524 )) ) + ( Xd_0__inst_mult_14_370  ) + ( Xd_0__inst_mult_14_369  ))
// Xd_0__inst_mult_14_373  = CARRY(( !Xd_0__inst_mult_14_516  $ (!Xd_0__inst_mult_14_520  $ (Xd_0__inst_mult_14_524 )) ) + ( Xd_0__inst_mult_14_370  ) + ( Xd_0__inst_mult_14_369  ))
// Xd_0__inst_mult_14_374  = SHARE((!Xd_0__inst_mult_14_516  & (Xd_0__inst_mult_14_520  & Xd_0__inst_mult_14_524 )) # (Xd_0__inst_mult_14_516  & ((Xd_0__inst_mult_14_524 ) # (Xd_0__inst_mult_14_520 ))))

	.dataa(!Xd_0__inst_mult_14_516 ),
	.datab(!Xd_0__inst_mult_14_520 ),
	.datac(!Xd_0__inst_mult_14_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_369 ),
	.sharein(Xd_0__inst_mult_14_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_372 ),
	.cout(Xd_0__inst_mult_14_373 ),
	.shareout(Xd_0__inst_mult_14_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_120 (
// Equation(s):
// Xd_0__inst_mult_15_380  = SUM(( !Xd_0__inst_mult_15_544  $ (!Xd_0__inst_mult_15_412  $ (Xd_0__inst_mult_15_548 )) ) + ( Xd_0__inst_mult_15_378  ) + ( Xd_0__inst_mult_15_377  ))
// Xd_0__inst_mult_15_381  = CARRY(( !Xd_0__inst_mult_15_544  $ (!Xd_0__inst_mult_15_412  $ (Xd_0__inst_mult_15_548 )) ) + ( Xd_0__inst_mult_15_378  ) + ( Xd_0__inst_mult_15_377  ))
// Xd_0__inst_mult_15_382  = SHARE((!Xd_0__inst_mult_15_544  & (Xd_0__inst_mult_15_412  & Xd_0__inst_mult_15_548 )) # (Xd_0__inst_mult_15_544  & ((Xd_0__inst_mult_15_548 ) # (Xd_0__inst_mult_15_412 ))))

	.dataa(!Xd_0__inst_mult_15_544 ),
	.datab(!Xd_0__inst_mult_15_412 ),
	.datac(!Xd_0__inst_mult_15_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_377 ),
	.sharein(Xd_0__inst_mult_15_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_380 ),
	.cout(Xd_0__inst_mult_15_381 ),
	.shareout(Xd_0__inst_mult_15_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_110 (
// Equation(s):
// Xd_0__inst_mult_10_352  = SUM(( !Xd_0__inst_mult_10_512  $ (!Xd_0__inst_mult_10_516  $ (Xd_0__inst_mult_10_520 )) ) + ( Xd_0__inst_mult_10_350  ) + ( Xd_0__inst_mult_10_349  ))
// Xd_0__inst_mult_10_353  = CARRY(( !Xd_0__inst_mult_10_512  $ (!Xd_0__inst_mult_10_516  $ (Xd_0__inst_mult_10_520 )) ) + ( Xd_0__inst_mult_10_350  ) + ( Xd_0__inst_mult_10_349  ))
// Xd_0__inst_mult_10_354  = SHARE((!Xd_0__inst_mult_10_512  & (Xd_0__inst_mult_10_516  & Xd_0__inst_mult_10_520 )) # (Xd_0__inst_mult_10_512  & ((Xd_0__inst_mult_10_520 ) # (Xd_0__inst_mult_10_516 ))))

	.dataa(!Xd_0__inst_mult_10_512 ),
	.datab(!Xd_0__inst_mult_10_516 ),
	.datac(!Xd_0__inst_mult_10_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_349 ),
	.sharein(Xd_0__inst_mult_10_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_352 ),
	.cout(Xd_0__inst_mult_10_353 ),
	.shareout(Xd_0__inst_mult_10_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_114 (
// Equation(s):
// Xd_0__inst_mult_11_356  = SUM(( !Xd_0__inst_mult_11_516  $ (!Xd_0__inst_mult_11_520  $ (Xd_0__inst_mult_11_524 )) ) + ( Xd_0__inst_mult_11_354  ) + ( Xd_0__inst_mult_11_353  ))
// Xd_0__inst_mult_11_357  = CARRY(( !Xd_0__inst_mult_11_516  $ (!Xd_0__inst_mult_11_520  $ (Xd_0__inst_mult_11_524 )) ) + ( Xd_0__inst_mult_11_354  ) + ( Xd_0__inst_mult_11_353  ))
// Xd_0__inst_mult_11_358  = SHARE((!Xd_0__inst_mult_11_516  & (Xd_0__inst_mult_11_520  & Xd_0__inst_mult_11_524 )) # (Xd_0__inst_mult_11_516  & ((Xd_0__inst_mult_11_524 ) # (Xd_0__inst_mult_11_520 ))))

	.dataa(!Xd_0__inst_mult_11_516 ),
	.datab(!Xd_0__inst_mult_11_520 ),
	.datac(!Xd_0__inst_mult_11_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_353 ),
	.sharein(Xd_0__inst_mult_11_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_356 ),
	.cout(Xd_0__inst_mult_11_357 ),
	.shareout(Xd_0__inst_mult_11_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_114 (
// Equation(s):
// Xd_0__inst_mult_8_356  = SUM(( !Xd_0__inst_mult_8_516  $ (!Xd_0__inst_mult_8_520  $ (Xd_0__inst_mult_8_524 )) ) + ( Xd_0__inst_mult_8_354  ) + ( Xd_0__inst_mult_8_353  ))
// Xd_0__inst_mult_8_357  = CARRY(( !Xd_0__inst_mult_8_516  $ (!Xd_0__inst_mult_8_520  $ (Xd_0__inst_mult_8_524 )) ) + ( Xd_0__inst_mult_8_354  ) + ( Xd_0__inst_mult_8_353  ))
// Xd_0__inst_mult_8_358  = SHARE((!Xd_0__inst_mult_8_516  & (Xd_0__inst_mult_8_520  & Xd_0__inst_mult_8_524 )) # (Xd_0__inst_mult_8_516  & ((Xd_0__inst_mult_8_524 ) # (Xd_0__inst_mult_8_520 ))))

	.dataa(!Xd_0__inst_mult_8_516 ),
	.datab(!Xd_0__inst_mult_8_520 ),
	.datac(!Xd_0__inst_mult_8_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_353 ),
	.sharein(Xd_0__inst_mult_8_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_356 ),
	.cout(Xd_0__inst_mult_8_357 ),
	.shareout(Xd_0__inst_mult_8_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_110 (
// Equation(s):
// Xd_0__inst_mult_9_352  = SUM(( !Xd_0__inst_mult_9_512  $ (!Xd_0__inst_mult_9_516  $ (Xd_0__inst_mult_9_520 )) ) + ( Xd_0__inst_mult_9_350  ) + ( Xd_0__inst_mult_9_349  ))
// Xd_0__inst_mult_9_353  = CARRY(( !Xd_0__inst_mult_9_512  $ (!Xd_0__inst_mult_9_516  $ (Xd_0__inst_mult_9_520 )) ) + ( Xd_0__inst_mult_9_350  ) + ( Xd_0__inst_mult_9_349  ))
// Xd_0__inst_mult_9_354  = SHARE((!Xd_0__inst_mult_9_512  & (Xd_0__inst_mult_9_516  & Xd_0__inst_mult_9_520 )) # (Xd_0__inst_mult_9_512  & ((Xd_0__inst_mult_9_520 ) # (Xd_0__inst_mult_9_516 ))))

	.dataa(!Xd_0__inst_mult_9_512 ),
	.datab(!Xd_0__inst_mult_9_516 ),
	.datac(!Xd_0__inst_mult_9_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_349 ),
	.sharein(Xd_0__inst_mult_9_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_352 ),
	.cout(Xd_0__inst_mult_9_353 ),
	.shareout(Xd_0__inst_mult_9_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_110 (
// Equation(s):
// Xd_0__inst_mult_6_352  = SUM(( !Xd_0__inst_mult_6_512  $ (!Xd_0__inst_mult_6_516  $ (Xd_0__inst_mult_6_520 )) ) + ( Xd_0__inst_mult_6_350  ) + ( Xd_0__inst_mult_6_349  ))
// Xd_0__inst_mult_6_353  = CARRY(( !Xd_0__inst_mult_6_512  $ (!Xd_0__inst_mult_6_516  $ (Xd_0__inst_mult_6_520 )) ) + ( Xd_0__inst_mult_6_350  ) + ( Xd_0__inst_mult_6_349  ))
// Xd_0__inst_mult_6_354  = SHARE((!Xd_0__inst_mult_6_512  & (Xd_0__inst_mult_6_516  & Xd_0__inst_mult_6_520 )) # (Xd_0__inst_mult_6_512  & ((Xd_0__inst_mult_6_520 ) # (Xd_0__inst_mult_6_516 ))))

	.dataa(!Xd_0__inst_mult_6_512 ),
	.datab(!Xd_0__inst_mult_6_516 ),
	.datac(!Xd_0__inst_mult_6_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_349 ),
	.sharein(Xd_0__inst_mult_6_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_352 ),
	.cout(Xd_0__inst_mult_6_353 ),
	.shareout(Xd_0__inst_mult_6_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_105 (
// Equation(s):
// Xd_0__inst_mult_7_332  = SUM(( !Xd_0__inst_mult_7_504  $ (((!din_b[87]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_326  ) + ( Xd_0__inst_mult_7_325  ))
// Xd_0__inst_mult_7_333  = CARRY(( !Xd_0__inst_mult_7_504  $ (((!din_b[87]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_326  ) + ( Xd_0__inst_mult_7_325  ))
// Xd_0__inst_mult_7_334  = SHARE((din_b[87] & (din_a[94] & Xd_0__inst_mult_7_504 )))

	.dataa(!din_b[87]),
	.datab(!din_a[94]),
	.datac(!Xd_0__inst_mult_7_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_325 ),
	.sharein(Xd_0__inst_mult_7_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_332 ),
	.cout(Xd_0__inst_mult_7_333 ),
	.shareout(Xd_0__inst_mult_7_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_106 (
// Equation(s):
// Xd_0__inst_mult_7_336  = SUM(( !Xd_0__inst_mult_7_508  $ (!Xd_0__inst_mult_7_512  $ (Xd_0__inst_mult_7_516 )) ) + ( Xd_0__inst_mult_7_330  ) + ( Xd_0__inst_mult_7_329  ))
// Xd_0__inst_mult_7_337  = CARRY(( !Xd_0__inst_mult_7_508  $ (!Xd_0__inst_mult_7_512  $ (Xd_0__inst_mult_7_516 )) ) + ( Xd_0__inst_mult_7_330  ) + ( Xd_0__inst_mult_7_329  ))
// Xd_0__inst_mult_7_338  = SHARE((!Xd_0__inst_mult_7_508  & (Xd_0__inst_mult_7_512  & Xd_0__inst_mult_7_516 )) # (Xd_0__inst_mult_7_508  & ((Xd_0__inst_mult_7_516 ) # (Xd_0__inst_mult_7_512 ))))

	.dataa(!Xd_0__inst_mult_7_508 ),
	.datab(!Xd_0__inst_mult_7_512 ),
	.datac(!Xd_0__inst_mult_7_516 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_329 ),
	.sharein(Xd_0__inst_mult_7_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_336 ),
	.cout(Xd_0__inst_mult_7_337 ),
	.shareout(Xd_0__inst_mult_7_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_117 (
// Equation(s):
// Xd_0__inst_mult_4_368  = SUM(( !Xd_0__inst_mult_4_536  $ (((!din_b[51]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_362  ) + ( Xd_0__inst_mult_4_361  ))
// Xd_0__inst_mult_4_369  = CARRY(( !Xd_0__inst_mult_4_536  $ (((!din_b[51]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_362  ) + ( Xd_0__inst_mult_4_361  ))
// Xd_0__inst_mult_4_370  = SHARE((din_b[51] & (din_a[58] & Xd_0__inst_mult_4_536 )))

	.dataa(!din_b[51]),
	.datab(!din_a[58]),
	.datac(!Xd_0__inst_mult_4_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_361 ),
	.sharein(Xd_0__inst_mult_4_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_368 ),
	.cout(Xd_0__inst_mult_4_369 ),
	.shareout(Xd_0__inst_mult_4_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_118 (
// Equation(s):
// Xd_0__inst_mult_4_372  = SUM(( !Xd_0__inst_mult_4_540  $ (!Xd_0__inst_mult_4_268  $ (Xd_0__inst_mult_4_544 )) ) + ( Xd_0__inst_mult_4_366  ) + ( Xd_0__inst_mult_4_365  ))
// Xd_0__inst_mult_4_373  = CARRY(( !Xd_0__inst_mult_4_540  $ (!Xd_0__inst_mult_4_268  $ (Xd_0__inst_mult_4_544 )) ) + ( Xd_0__inst_mult_4_366  ) + ( Xd_0__inst_mult_4_365  ))
// Xd_0__inst_mult_4_374  = SHARE((!Xd_0__inst_mult_4_540  & (Xd_0__inst_mult_4_268  & Xd_0__inst_mult_4_544 )) # (Xd_0__inst_mult_4_540  & ((Xd_0__inst_mult_4_544 ) # (Xd_0__inst_mult_4_268 ))))

	.dataa(!Xd_0__inst_mult_4_540 ),
	.datab(!Xd_0__inst_mult_4_268 ),
	.datac(!Xd_0__inst_mult_4_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_365 ),
	.sharein(Xd_0__inst_mult_4_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_372 ),
	.cout(Xd_0__inst_mult_4_373 ),
	.shareout(Xd_0__inst_mult_4_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_105 (
// Equation(s):
// Xd_0__inst_mult_5_332  = SUM(( !Xd_0__inst_mult_5_504  $ (((!din_b[63]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_326  ) + ( Xd_0__inst_mult_5_325  ))
// Xd_0__inst_mult_5_333  = CARRY(( !Xd_0__inst_mult_5_504  $ (((!din_b[63]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_326  ) + ( Xd_0__inst_mult_5_325  ))
// Xd_0__inst_mult_5_334  = SHARE((din_b[63] & (din_a[70] & Xd_0__inst_mult_5_504 )))

	.dataa(!din_b[63]),
	.datab(!din_a[70]),
	.datac(!Xd_0__inst_mult_5_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_325 ),
	.sharein(Xd_0__inst_mult_5_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_332 ),
	.cout(Xd_0__inst_mult_5_333 ),
	.shareout(Xd_0__inst_mult_5_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_106 (
// Equation(s):
// Xd_0__inst_mult_5_336  = SUM(( !Xd_0__inst_mult_5_508  $ (!Xd_0__inst_mult_5_512  $ (Xd_0__inst_mult_5_516 )) ) + ( Xd_0__inst_mult_5_330  ) + ( Xd_0__inst_mult_5_329  ))
// Xd_0__inst_mult_5_337  = CARRY(( !Xd_0__inst_mult_5_508  $ (!Xd_0__inst_mult_5_512  $ (Xd_0__inst_mult_5_516 )) ) + ( Xd_0__inst_mult_5_330  ) + ( Xd_0__inst_mult_5_329  ))
// Xd_0__inst_mult_5_338  = SHARE((!Xd_0__inst_mult_5_508  & (Xd_0__inst_mult_5_512  & Xd_0__inst_mult_5_516 )) # (Xd_0__inst_mult_5_508  & ((Xd_0__inst_mult_5_516 ) # (Xd_0__inst_mult_5_512 ))))

	.dataa(!Xd_0__inst_mult_5_508 ),
	.datab(!Xd_0__inst_mult_5_512 ),
	.datac(!Xd_0__inst_mult_5_516 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_329 ),
	.sharein(Xd_0__inst_mult_5_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_336 ),
	.cout(Xd_0__inst_mult_5_337 ),
	.shareout(Xd_0__inst_mult_5_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_109 (
// Equation(s):
// Xd_0__inst_mult_2_336  = SUM(( !Xd_0__inst_mult_2_508  $ (((!din_b[27]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_330  ) + ( Xd_0__inst_mult_2_329  ))
// Xd_0__inst_mult_2_337  = CARRY(( !Xd_0__inst_mult_2_508  $ (((!din_b[27]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_330  ) + ( Xd_0__inst_mult_2_329  ))
// Xd_0__inst_mult_2_338  = SHARE((din_b[27] & (din_a[34] & Xd_0__inst_mult_2_508 )))

	.dataa(!din_b[27]),
	.datab(!din_a[34]),
	.datac(!Xd_0__inst_mult_2_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_329 ),
	.sharein(Xd_0__inst_mult_2_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_336 ),
	.cout(Xd_0__inst_mult_2_337 ),
	.shareout(Xd_0__inst_mult_2_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_110 (
// Equation(s):
// Xd_0__inst_mult_2_340  = SUM(( !Xd_0__inst_mult_2_512  $ (!Xd_0__inst_mult_2_516  $ (Xd_0__inst_mult_2_520 )) ) + ( Xd_0__inst_mult_2_334  ) + ( Xd_0__inst_mult_2_333  ))
// Xd_0__inst_mult_2_341  = CARRY(( !Xd_0__inst_mult_2_512  $ (!Xd_0__inst_mult_2_516  $ (Xd_0__inst_mult_2_520 )) ) + ( Xd_0__inst_mult_2_334  ) + ( Xd_0__inst_mult_2_333  ))
// Xd_0__inst_mult_2_342  = SHARE((!Xd_0__inst_mult_2_512  & (Xd_0__inst_mult_2_516  & Xd_0__inst_mult_2_520 )) # (Xd_0__inst_mult_2_512  & ((Xd_0__inst_mult_2_520 ) # (Xd_0__inst_mult_2_516 ))))

	.dataa(!Xd_0__inst_mult_2_512 ),
	.datab(!Xd_0__inst_mult_2_516 ),
	.datac(!Xd_0__inst_mult_2_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_333 ),
	.sharein(Xd_0__inst_mult_2_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_340 ),
	.cout(Xd_0__inst_mult_2_341 ),
	.shareout(Xd_0__inst_mult_2_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_105 (
// Equation(s):
// Xd_0__inst_mult_3_332  = SUM(( !Xd_0__inst_mult_3_504  $ (((!din_b[39]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_326  ) + ( Xd_0__inst_mult_3_325  ))
// Xd_0__inst_mult_3_333  = CARRY(( !Xd_0__inst_mult_3_504  $ (((!din_b[39]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_326  ) + ( Xd_0__inst_mult_3_325  ))
// Xd_0__inst_mult_3_334  = SHARE((din_b[39] & (din_a[46] & Xd_0__inst_mult_3_504 )))

	.dataa(!din_b[39]),
	.datab(!din_a[46]),
	.datac(!Xd_0__inst_mult_3_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_325 ),
	.sharein(Xd_0__inst_mult_3_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_332 ),
	.cout(Xd_0__inst_mult_3_333 ),
	.shareout(Xd_0__inst_mult_3_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_106 (
// Equation(s):
// Xd_0__inst_mult_3_336  = SUM(( !Xd_0__inst_mult_3_508  $ (!Xd_0__inst_mult_3_512  $ (Xd_0__inst_mult_3_516 )) ) + ( Xd_0__inst_mult_3_330  ) + ( Xd_0__inst_mult_3_329  ))
// Xd_0__inst_mult_3_337  = CARRY(( !Xd_0__inst_mult_3_508  $ (!Xd_0__inst_mult_3_512  $ (Xd_0__inst_mult_3_516 )) ) + ( Xd_0__inst_mult_3_330  ) + ( Xd_0__inst_mult_3_329  ))
// Xd_0__inst_mult_3_338  = SHARE((!Xd_0__inst_mult_3_508  & (Xd_0__inst_mult_3_512  & Xd_0__inst_mult_3_516 )) # (Xd_0__inst_mult_3_508  & ((Xd_0__inst_mult_3_516 ) # (Xd_0__inst_mult_3_512 ))))

	.dataa(!Xd_0__inst_mult_3_508 ),
	.datab(!Xd_0__inst_mult_3_512 ),
	.datac(!Xd_0__inst_mult_3_516 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_329 ),
	.sharein(Xd_0__inst_mult_3_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_336 ),
	.cout(Xd_0__inst_mult_3_337 ),
	.shareout(Xd_0__inst_mult_3_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_109 (
// Equation(s):
// Xd_0__inst_mult_0_336  = SUM(( !Xd_0__inst_mult_0_508  $ (((!din_b[3]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_330  ) + ( Xd_0__inst_mult_0_329  ))
// Xd_0__inst_mult_0_337  = CARRY(( !Xd_0__inst_mult_0_508  $ (((!din_b[3]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_330  ) + ( Xd_0__inst_mult_0_329  ))
// Xd_0__inst_mult_0_338  = SHARE((din_b[3] & (din_a[10] & Xd_0__inst_mult_0_508 )))

	.dataa(!din_b[3]),
	.datab(!din_a[10]),
	.datac(!Xd_0__inst_mult_0_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_329 ),
	.sharein(Xd_0__inst_mult_0_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_336 ),
	.cout(Xd_0__inst_mult_0_337 ),
	.shareout(Xd_0__inst_mult_0_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_110 (
// Equation(s):
// Xd_0__inst_mult_0_340  = SUM(( !Xd_0__inst_mult_0_512  $ (!Xd_0__inst_mult_0_516  $ (Xd_0__inst_mult_0_520 )) ) + ( Xd_0__inst_mult_0_334  ) + ( Xd_0__inst_mult_0_333  ))
// Xd_0__inst_mult_0_341  = CARRY(( !Xd_0__inst_mult_0_512  $ (!Xd_0__inst_mult_0_516  $ (Xd_0__inst_mult_0_520 )) ) + ( Xd_0__inst_mult_0_334  ) + ( Xd_0__inst_mult_0_333  ))
// Xd_0__inst_mult_0_342  = SHARE((!Xd_0__inst_mult_0_512  & (Xd_0__inst_mult_0_516  & Xd_0__inst_mult_0_520 )) # (Xd_0__inst_mult_0_512  & ((Xd_0__inst_mult_0_520 ) # (Xd_0__inst_mult_0_516 ))))

	.dataa(!Xd_0__inst_mult_0_512 ),
	.datab(!Xd_0__inst_mult_0_516 ),
	.datac(!Xd_0__inst_mult_0_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_333 ),
	.sharein(Xd_0__inst_mult_0_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_340 ),
	.cout(Xd_0__inst_mult_0_341 ),
	.shareout(Xd_0__inst_mult_0_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_109 (
// Equation(s):
// Xd_0__inst_mult_1_336  = SUM(( !Xd_0__inst_mult_1_508  $ (((!din_b[15]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_330  ) + ( Xd_0__inst_mult_1_329  ))
// Xd_0__inst_mult_1_337  = CARRY(( !Xd_0__inst_mult_1_508  $ (((!din_b[15]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_330  ) + ( Xd_0__inst_mult_1_329  ))
// Xd_0__inst_mult_1_338  = SHARE((din_b[15] & (din_a[22] & Xd_0__inst_mult_1_508 )))

	.dataa(!din_b[15]),
	.datab(!din_a[22]),
	.datac(!Xd_0__inst_mult_1_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_329 ),
	.sharein(Xd_0__inst_mult_1_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_336 ),
	.cout(Xd_0__inst_mult_1_337 ),
	.shareout(Xd_0__inst_mult_1_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_110 (
// Equation(s):
// Xd_0__inst_mult_1_340  = SUM(( !Xd_0__inst_mult_1_512  $ (!Xd_0__inst_mult_1_516  $ (Xd_0__inst_mult_1_520 )) ) + ( Xd_0__inst_mult_1_334  ) + ( Xd_0__inst_mult_1_333  ))
// Xd_0__inst_mult_1_341  = CARRY(( !Xd_0__inst_mult_1_512  $ (!Xd_0__inst_mult_1_516  $ (Xd_0__inst_mult_1_520 )) ) + ( Xd_0__inst_mult_1_334  ) + ( Xd_0__inst_mult_1_333  ))
// Xd_0__inst_mult_1_342  = SHARE((!Xd_0__inst_mult_1_512  & (Xd_0__inst_mult_1_516  & Xd_0__inst_mult_1_520 )) # (Xd_0__inst_mult_1_512  & ((Xd_0__inst_mult_1_520 ) # (Xd_0__inst_mult_1_516 ))))

	.dataa(!Xd_0__inst_mult_1_512 ),
	.datab(!Xd_0__inst_mult_1_516 ),
	.datac(!Xd_0__inst_mult_1_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_333 ),
	.sharein(Xd_0__inst_mult_1_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_340 ),
	.cout(Xd_0__inst_mult_1_341 ),
	.shareout(Xd_0__inst_mult_1_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_117 (
// Equation(s):
// Xd_0__inst_mult_12_380  = SUM(( !Xd_0__inst_mult_12_548  $ (!Xd_0__inst_mult_12_300  $ (Xd_0__inst_mult_12_552 )) ) + ( Xd_0__inst_mult_12_378  ) + ( Xd_0__inst_mult_12_377  ))
// Xd_0__inst_mult_12_381  = CARRY(( !Xd_0__inst_mult_12_548  $ (!Xd_0__inst_mult_12_300  $ (Xd_0__inst_mult_12_552 )) ) + ( Xd_0__inst_mult_12_378  ) + ( Xd_0__inst_mult_12_377  ))
// Xd_0__inst_mult_12_382  = SHARE((!Xd_0__inst_mult_12_548  & (Xd_0__inst_mult_12_300  & Xd_0__inst_mult_12_552 )) # (Xd_0__inst_mult_12_548  & ((Xd_0__inst_mult_12_552 ) # (Xd_0__inst_mult_12_300 ))))

	.dataa(!Xd_0__inst_mult_12_548 ),
	.datab(!Xd_0__inst_mult_12_300 ),
	.datac(!Xd_0__inst_mult_12_552 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_377 ),
	.sharein(Xd_0__inst_mult_12_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_380 ),
	.cout(Xd_0__inst_mult_12_381 ),
	.shareout(Xd_0__inst_mult_12_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_115 (
// Equation(s):
// Xd_0__inst_mult_13_360  = SUM(( !Xd_0__inst_mult_13_528  $ (!Xd_0__inst_mult_13_532  $ (Xd_0__inst_mult_13_536 )) ) + ( Xd_0__inst_mult_13_358  ) + ( Xd_0__inst_mult_13_357  ))
// Xd_0__inst_mult_13_361  = CARRY(( !Xd_0__inst_mult_13_528  $ (!Xd_0__inst_mult_13_532  $ (Xd_0__inst_mult_13_536 )) ) + ( Xd_0__inst_mult_13_358  ) + ( Xd_0__inst_mult_13_357  ))
// Xd_0__inst_mult_13_362  = SHARE((!Xd_0__inst_mult_13_528  & (Xd_0__inst_mult_13_532  & Xd_0__inst_mult_13_536 )) # (Xd_0__inst_mult_13_528  & ((Xd_0__inst_mult_13_536 ) # (Xd_0__inst_mult_13_532 ))))

	.dataa(!Xd_0__inst_mult_13_528 ),
	.datab(!Xd_0__inst_mult_13_532 ),
	.datac(!Xd_0__inst_mult_13_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_357 ),
	.sharein(Xd_0__inst_mult_13_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_360 ),
	.cout(Xd_0__inst_mult_13_361 ),
	.shareout(Xd_0__inst_mult_13_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_119 (
// Equation(s):
// Xd_0__inst_mult_14_376  = SUM(( !Xd_0__inst_mult_14_528  $ (!Xd_0__inst_mult_14_532  $ (Xd_0__inst_mult_14_536 )) ) + ( Xd_0__inst_mult_14_374  ) + ( Xd_0__inst_mult_14_373  ))
// Xd_0__inst_mult_14_377  = CARRY(( !Xd_0__inst_mult_14_528  $ (!Xd_0__inst_mult_14_532  $ (Xd_0__inst_mult_14_536 )) ) + ( Xd_0__inst_mult_14_374  ) + ( Xd_0__inst_mult_14_373  ))
// Xd_0__inst_mult_14_378  = SHARE((!Xd_0__inst_mult_14_528  & (Xd_0__inst_mult_14_532  & Xd_0__inst_mult_14_536 )) # (Xd_0__inst_mult_14_528  & ((Xd_0__inst_mult_14_536 ) # (Xd_0__inst_mult_14_532 ))))

	.dataa(!Xd_0__inst_mult_14_528 ),
	.datab(!Xd_0__inst_mult_14_532 ),
	.datac(!Xd_0__inst_mult_14_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_373 ),
	.sharein(Xd_0__inst_mult_14_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_376 ),
	.cout(Xd_0__inst_mult_14_377 ),
	.shareout(Xd_0__inst_mult_14_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_121 (
// Equation(s):
// Xd_0__inst_mult_15_384  = SUM(( !Xd_0__inst_mult_15_552  $ (!Xd_0__inst_mult_15_296  $ (Xd_0__inst_mult_15_556 )) ) + ( Xd_0__inst_mult_15_382  ) + ( Xd_0__inst_mult_15_381  ))
// Xd_0__inst_mult_15_385  = CARRY(( !Xd_0__inst_mult_15_552  $ (!Xd_0__inst_mult_15_296  $ (Xd_0__inst_mult_15_556 )) ) + ( Xd_0__inst_mult_15_382  ) + ( Xd_0__inst_mult_15_381  ))
// Xd_0__inst_mult_15_386  = SHARE((!Xd_0__inst_mult_15_552  & (Xd_0__inst_mult_15_296  & Xd_0__inst_mult_15_556 )) # (Xd_0__inst_mult_15_552  & ((Xd_0__inst_mult_15_556 ) # (Xd_0__inst_mult_15_296 ))))

	.dataa(!Xd_0__inst_mult_15_552 ),
	.datab(!Xd_0__inst_mult_15_296 ),
	.datac(!Xd_0__inst_mult_15_556 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_381 ),
	.sharein(Xd_0__inst_mult_15_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_384 ),
	.cout(Xd_0__inst_mult_15_385 ),
	.shareout(Xd_0__inst_mult_15_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_111 (
// Equation(s):
// Xd_0__inst_mult_10_356  = SUM(( !Xd_0__inst_mult_10_524  $ (!Xd_0__inst_mult_10_528  $ (Xd_0__inst_mult_10_532 )) ) + ( Xd_0__inst_mult_10_354  ) + ( Xd_0__inst_mult_10_353  ))
// Xd_0__inst_mult_10_357  = CARRY(( !Xd_0__inst_mult_10_524  $ (!Xd_0__inst_mult_10_528  $ (Xd_0__inst_mult_10_532 )) ) + ( Xd_0__inst_mult_10_354  ) + ( Xd_0__inst_mult_10_353  ))
// Xd_0__inst_mult_10_358  = SHARE((!Xd_0__inst_mult_10_524  & (Xd_0__inst_mult_10_528  & Xd_0__inst_mult_10_532 )) # (Xd_0__inst_mult_10_524  & ((Xd_0__inst_mult_10_532 ) # (Xd_0__inst_mult_10_528 ))))

	.dataa(!Xd_0__inst_mult_10_524 ),
	.datab(!Xd_0__inst_mult_10_528 ),
	.datac(!Xd_0__inst_mult_10_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_353 ),
	.sharein(Xd_0__inst_mult_10_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_356 ),
	.cout(Xd_0__inst_mult_10_357 ),
	.shareout(Xd_0__inst_mult_10_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_115 (
// Equation(s):
// Xd_0__inst_mult_11_360  = SUM(( !Xd_0__inst_mult_11_528  $ (!Xd_0__inst_mult_11_532  $ (Xd_0__inst_mult_11_536 )) ) + ( Xd_0__inst_mult_11_358  ) + ( Xd_0__inst_mult_11_357  ))
// Xd_0__inst_mult_11_361  = CARRY(( !Xd_0__inst_mult_11_528  $ (!Xd_0__inst_mult_11_532  $ (Xd_0__inst_mult_11_536 )) ) + ( Xd_0__inst_mult_11_358  ) + ( Xd_0__inst_mult_11_357  ))
// Xd_0__inst_mult_11_362  = SHARE((!Xd_0__inst_mult_11_528  & (Xd_0__inst_mult_11_532  & Xd_0__inst_mult_11_536 )) # (Xd_0__inst_mult_11_528  & ((Xd_0__inst_mult_11_536 ) # (Xd_0__inst_mult_11_532 ))))

	.dataa(!Xd_0__inst_mult_11_528 ),
	.datab(!Xd_0__inst_mult_11_532 ),
	.datac(!Xd_0__inst_mult_11_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_357 ),
	.sharein(Xd_0__inst_mult_11_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_360 ),
	.cout(Xd_0__inst_mult_11_361 ),
	.shareout(Xd_0__inst_mult_11_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_115 (
// Equation(s):
// Xd_0__inst_mult_8_360  = SUM(( !Xd_0__inst_mult_8_528  $ (!Xd_0__inst_mult_8_532  $ (Xd_0__inst_mult_8_536 )) ) + ( Xd_0__inst_mult_8_358  ) + ( Xd_0__inst_mult_8_357  ))
// Xd_0__inst_mult_8_361  = CARRY(( !Xd_0__inst_mult_8_528  $ (!Xd_0__inst_mult_8_532  $ (Xd_0__inst_mult_8_536 )) ) + ( Xd_0__inst_mult_8_358  ) + ( Xd_0__inst_mult_8_357  ))
// Xd_0__inst_mult_8_362  = SHARE((!Xd_0__inst_mult_8_528  & (Xd_0__inst_mult_8_532  & Xd_0__inst_mult_8_536 )) # (Xd_0__inst_mult_8_528  & ((Xd_0__inst_mult_8_536 ) # (Xd_0__inst_mult_8_532 ))))

	.dataa(!Xd_0__inst_mult_8_528 ),
	.datab(!Xd_0__inst_mult_8_532 ),
	.datac(!Xd_0__inst_mult_8_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_357 ),
	.sharein(Xd_0__inst_mult_8_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_360 ),
	.cout(Xd_0__inst_mult_8_361 ),
	.shareout(Xd_0__inst_mult_8_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_111 (
// Equation(s):
// Xd_0__inst_mult_9_356  = SUM(( !Xd_0__inst_mult_9_524  $ (!Xd_0__inst_mult_9_528  $ (Xd_0__inst_mult_9_532 )) ) + ( Xd_0__inst_mult_9_354  ) + ( Xd_0__inst_mult_9_353  ))
// Xd_0__inst_mult_9_357  = CARRY(( !Xd_0__inst_mult_9_524  $ (!Xd_0__inst_mult_9_528  $ (Xd_0__inst_mult_9_532 )) ) + ( Xd_0__inst_mult_9_354  ) + ( Xd_0__inst_mult_9_353  ))
// Xd_0__inst_mult_9_358  = SHARE((!Xd_0__inst_mult_9_524  & (Xd_0__inst_mult_9_528  & Xd_0__inst_mult_9_532 )) # (Xd_0__inst_mult_9_524  & ((Xd_0__inst_mult_9_532 ) # (Xd_0__inst_mult_9_528 ))))

	.dataa(!Xd_0__inst_mult_9_524 ),
	.datab(!Xd_0__inst_mult_9_528 ),
	.datac(!Xd_0__inst_mult_9_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_353 ),
	.sharein(Xd_0__inst_mult_9_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_356 ),
	.cout(Xd_0__inst_mult_9_357 ),
	.shareout(Xd_0__inst_mult_9_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_111 (
// Equation(s):
// Xd_0__inst_mult_6_356  = SUM(( !Xd_0__inst_mult_6_524  $ (!Xd_0__inst_mult_6_528  $ (Xd_0__inst_mult_6_532 )) ) + ( Xd_0__inst_mult_6_354  ) + ( Xd_0__inst_mult_6_353  ))
// Xd_0__inst_mult_6_357  = CARRY(( !Xd_0__inst_mult_6_524  $ (!Xd_0__inst_mult_6_528  $ (Xd_0__inst_mult_6_532 )) ) + ( Xd_0__inst_mult_6_354  ) + ( Xd_0__inst_mult_6_353  ))
// Xd_0__inst_mult_6_358  = SHARE((!Xd_0__inst_mult_6_524  & (Xd_0__inst_mult_6_528  & Xd_0__inst_mult_6_532 )) # (Xd_0__inst_mult_6_524  & ((Xd_0__inst_mult_6_532 ) # (Xd_0__inst_mult_6_528 ))))

	.dataa(!Xd_0__inst_mult_6_524 ),
	.datab(!Xd_0__inst_mult_6_528 ),
	.datac(!Xd_0__inst_mult_6_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_353 ),
	.sharein(Xd_0__inst_mult_6_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_356 ),
	.cout(Xd_0__inst_mult_6_357 ),
	.shareout(Xd_0__inst_mult_6_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_107 (
// Equation(s):
// Xd_0__inst_mult_7_340  = SUM(( !Xd_0__inst_mult_7_520  $ (((!din_b[88]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_334  ) + ( Xd_0__inst_mult_7_333  ))
// Xd_0__inst_mult_7_341  = CARRY(( !Xd_0__inst_mult_7_520  $ (((!din_b[88]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_334  ) + ( Xd_0__inst_mult_7_333  ))
// Xd_0__inst_mult_7_342  = SHARE((din_b[88] & (din_a[94] & Xd_0__inst_mult_7_520 )))

	.dataa(!din_b[88]),
	.datab(!din_a[94]),
	.datac(!Xd_0__inst_mult_7_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_333 ),
	.sharein(Xd_0__inst_mult_7_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_340 ),
	.cout(Xd_0__inst_mult_7_341 ),
	.shareout(Xd_0__inst_mult_7_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_108 (
// Equation(s):
// Xd_0__inst_mult_7_344  = SUM(( !Xd_0__inst_mult_7_524  $ (!Xd_0__inst_mult_7_528  $ (Xd_0__inst_mult_7_532 )) ) + ( Xd_0__inst_mult_7_338  ) + ( Xd_0__inst_mult_7_337  ))
// Xd_0__inst_mult_7_345  = CARRY(( !Xd_0__inst_mult_7_524  $ (!Xd_0__inst_mult_7_528  $ (Xd_0__inst_mult_7_532 )) ) + ( Xd_0__inst_mult_7_338  ) + ( Xd_0__inst_mult_7_337  ))
// Xd_0__inst_mult_7_346  = SHARE((!Xd_0__inst_mult_7_524  & (Xd_0__inst_mult_7_528  & Xd_0__inst_mult_7_532 )) # (Xd_0__inst_mult_7_524  & ((Xd_0__inst_mult_7_532 ) # (Xd_0__inst_mult_7_528 ))))

	.dataa(!Xd_0__inst_mult_7_524 ),
	.datab(!Xd_0__inst_mult_7_528 ),
	.datac(!Xd_0__inst_mult_7_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_337 ),
	.sharein(Xd_0__inst_mult_7_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_344 ),
	.cout(Xd_0__inst_mult_7_345 ),
	.shareout(Xd_0__inst_mult_7_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_119 (
// Equation(s):
// Xd_0__inst_mult_4_376  = SUM(( !Xd_0__inst_mult_4_548  $ (((!din_b[52]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_370  ) + ( Xd_0__inst_mult_4_369  ))
// Xd_0__inst_mult_4_377  = CARRY(( !Xd_0__inst_mult_4_548  $ (((!din_b[52]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_370  ) + ( Xd_0__inst_mult_4_369  ))
// Xd_0__inst_mult_4_378  = SHARE((din_b[52] & (din_a[58] & Xd_0__inst_mult_4_548 )))

	.dataa(!din_b[52]),
	.datab(!din_a[58]),
	.datac(!Xd_0__inst_mult_4_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_369 ),
	.sharein(Xd_0__inst_mult_4_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_376 ),
	.cout(Xd_0__inst_mult_4_377 ),
	.shareout(Xd_0__inst_mult_4_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_120 (
// Equation(s):
// Xd_0__inst_mult_4_380  = SUM(( !Xd_0__inst_mult_4_552  $ (!Xd_0__inst_mult_4_192  $ (Xd_0__inst_mult_4_556 )) ) + ( Xd_0__inst_mult_4_374  ) + ( Xd_0__inst_mult_4_373  ))
// Xd_0__inst_mult_4_381  = CARRY(( !Xd_0__inst_mult_4_552  $ (!Xd_0__inst_mult_4_192  $ (Xd_0__inst_mult_4_556 )) ) + ( Xd_0__inst_mult_4_374  ) + ( Xd_0__inst_mult_4_373  ))
// Xd_0__inst_mult_4_382  = SHARE((!Xd_0__inst_mult_4_552  & (Xd_0__inst_mult_4_192  & Xd_0__inst_mult_4_556 )) # (Xd_0__inst_mult_4_552  & ((Xd_0__inst_mult_4_556 ) # (Xd_0__inst_mult_4_192 ))))

	.dataa(!Xd_0__inst_mult_4_552 ),
	.datab(!Xd_0__inst_mult_4_192 ),
	.datac(!Xd_0__inst_mult_4_556 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_373 ),
	.sharein(Xd_0__inst_mult_4_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_380 ),
	.cout(Xd_0__inst_mult_4_381 ),
	.shareout(Xd_0__inst_mult_4_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_107 (
// Equation(s):
// Xd_0__inst_mult_5_340  = SUM(( !Xd_0__inst_mult_5_520  $ (((!din_b[64]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_334  ) + ( Xd_0__inst_mult_5_333  ))
// Xd_0__inst_mult_5_341  = CARRY(( !Xd_0__inst_mult_5_520  $ (((!din_b[64]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_334  ) + ( Xd_0__inst_mult_5_333  ))
// Xd_0__inst_mult_5_342  = SHARE((din_b[64] & (din_a[70] & Xd_0__inst_mult_5_520 )))

	.dataa(!din_b[64]),
	.datab(!din_a[70]),
	.datac(!Xd_0__inst_mult_5_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_333 ),
	.sharein(Xd_0__inst_mult_5_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_340 ),
	.cout(Xd_0__inst_mult_5_341 ),
	.shareout(Xd_0__inst_mult_5_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_108 (
// Equation(s):
// Xd_0__inst_mult_5_344  = SUM(( !Xd_0__inst_mult_5_524  $ (!Xd_0__inst_mult_5_528  $ (Xd_0__inst_mult_5_532 )) ) + ( Xd_0__inst_mult_5_338  ) + ( Xd_0__inst_mult_5_337  ))
// Xd_0__inst_mult_5_345  = CARRY(( !Xd_0__inst_mult_5_524  $ (!Xd_0__inst_mult_5_528  $ (Xd_0__inst_mult_5_532 )) ) + ( Xd_0__inst_mult_5_338  ) + ( Xd_0__inst_mult_5_337  ))
// Xd_0__inst_mult_5_346  = SHARE((!Xd_0__inst_mult_5_524  & (Xd_0__inst_mult_5_528  & Xd_0__inst_mult_5_532 )) # (Xd_0__inst_mult_5_524  & ((Xd_0__inst_mult_5_532 ) # (Xd_0__inst_mult_5_528 ))))

	.dataa(!Xd_0__inst_mult_5_524 ),
	.datab(!Xd_0__inst_mult_5_528 ),
	.datac(!Xd_0__inst_mult_5_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_337 ),
	.sharein(Xd_0__inst_mult_5_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_344 ),
	.cout(Xd_0__inst_mult_5_345 ),
	.shareout(Xd_0__inst_mult_5_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_111 (
// Equation(s):
// Xd_0__inst_mult_2_344  = SUM(( !Xd_0__inst_mult_2_524  $ (((!din_b[28]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_338  ) + ( Xd_0__inst_mult_2_337  ))
// Xd_0__inst_mult_2_345  = CARRY(( !Xd_0__inst_mult_2_524  $ (((!din_b[28]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_338  ) + ( Xd_0__inst_mult_2_337  ))
// Xd_0__inst_mult_2_346  = SHARE((din_b[28] & (din_a[34] & Xd_0__inst_mult_2_524 )))

	.dataa(!din_b[28]),
	.datab(!din_a[34]),
	.datac(!Xd_0__inst_mult_2_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_337 ),
	.sharein(Xd_0__inst_mult_2_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_344 ),
	.cout(Xd_0__inst_mult_2_345 ),
	.shareout(Xd_0__inst_mult_2_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_112 (
// Equation(s):
// Xd_0__inst_mult_2_348  = SUM(( !Xd_0__inst_mult_2_528  $ (!Xd_0__inst_mult_2_532  $ (Xd_0__inst_mult_2_536 )) ) + ( Xd_0__inst_mult_2_342  ) + ( Xd_0__inst_mult_2_341  ))
// Xd_0__inst_mult_2_349  = CARRY(( !Xd_0__inst_mult_2_528  $ (!Xd_0__inst_mult_2_532  $ (Xd_0__inst_mult_2_536 )) ) + ( Xd_0__inst_mult_2_342  ) + ( Xd_0__inst_mult_2_341  ))
// Xd_0__inst_mult_2_350  = SHARE((!Xd_0__inst_mult_2_528  & (Xd_0__inst_mult_2_532  & Xd_0__inst_mult_2_536 )) # (Xd_0__inst_mult_2_528  & ((Xd_0__inst_mult_2_536 ) # (Xd_0__inst_mult_2_532 ))))

	.dataa(!Xd_0__inst_mult_2_528 ),
	.datab(!Xd_0__inst_mult_2_532 ),
	.datac(!Xd_0__inst_mult_2_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_341 ),
	.sharein(Xd_0__inst_mult_2_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_348 ),
	.cout(Xd_0__inst_mult_2_349 ),
	.shareout(Xd_0__inst_mult_2_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_107 (
// Equation(s):
// Xd_0__inst_mult_3_340  = SUM(( !Xd_0__inst_mult_3_520  $ (((!din_b[40]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_334  ) + ( Xd_0__inst_mult_3_333  ))
// Xd_0__inst_mult_3_341  = CARRY(( !Xd_0__inst_mult_3_520  $ (((!din_b[40]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_334  ) + ( Xd_0__inst_mult_3_333  ))
// Xd_0__inst_mult_3_342  = SHARE((din_b[40] & (din_a[46] & Xd_0__inst_mult_3_520 )))

	.dataa(!din_b[40]),
	.datab(!din_a[46]),
	.datac(!Xd_0__inst_mult_3_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_333 ),
	.sharein(Xd_0__inst_mult_3_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_340 ),
	.cout(Xd_0__inst_mult_3_341 ),
	.shareout(Xd_0__inst_mult_3_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_108 (
// Equation(s):
// Xd_0__inst_mult_3_344  = SUM(( !Xd_0__inst_mult_3_524  $ (!Xd_0__inst_mult_3_528  $ (Xd_0__inst_mult_3_532 )) ) + ( Xd_0__inst_mult_3_338  ) + ( Xd_0__inst_mult_3_337  ))
// Xd_0__inst_mult_3_345  = CARRY(( !Xd_0__inst_mult_3_524  $ (!Xd_0__inst_mult_3_528  $ (Xd_0__inst_mult_3_532 )) ) + ( Xd_0__inst_mult_3_338  ) + ( Xd_0__inst_mult_3_337  ))
// Xd_0__inst_mult_3_346  = SHARE((!Xd_0__inst_mult_3_524  & (Xd_0__inst_mult_3_528  & Xd_0__inst_mult_3_532 )) # (Xd_0__inst_mult_3_524  & ((Xd_0__inst_mult_3_532 ) # (Xd_0__inst_mult_3_528 ))))

	.dataa(!Xd_0__inst_mult_3_524 ),
	.datab(!Xd_0__inst_mult_3_528 ),
	.datac(!Xd_0__inst_mult_3_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_337 ),
	.sharein(Xd_0__inst_mult_3_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_344 ),
	.cout(Xd_0__inst_mult_3_345 ),
	.shareout(Xd_0__inst_mult_3_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_111 (
// Equation(s):
// Xd_0__inst_mult_0_344  = SUM(( !Xd_0__inst_mult_0_524  $ (((!din_b[4]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_338  ) + ( Xd_0__inst_mult_0_337  ))
// Xd_0__inst_mult_0_345  = CARRY(( !Xd_0__inst_mult_0_524  $ (((!din_b[4]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_338  ) + ( Xd_0__inst_mult_0_337  ))
// Xd_0__inst_mult_0_346  = SHARE((din_b[4] & (din_a[10] & Xd_0__inst_mult_0_524 )))

	.dataa(!din_b[4]),
	.datab(!din_a[10]),
	.datac(!Xd_0__inst_mult_0_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_337 ),
	.sharein(Xd_0__inst_mult_0_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_344 ),
	.cout(Xd_0__inst_mult_0_345 ),
	.shareout(Xd_0__inst_mult_0_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_112 (
// Equation(s):
// Xd_0__inst_mult_0_348  = SUM(( !Xd_0__inst_mult_0_528  $ (!Xd_0__inst_mult_0_532  $ (Xd_0__inst_mult_0_536 )) ) + ( Xd_0__inst_mult_0_342  ) + ( Xd_0__inst_mult_0_341  ))
// Xd_0__inst_mult_0_349  = CARRY(( !Xd_0__inst_mult_0_528  $ (!Xd_0__inst_mult_0_532  $ (Xd_0__inst_mult_0_536 )) ) + ( Xd_0__inst_mult_0_342  ) + ( Xd_0__inst_mult_0_341  ))
// Xd_0__inst_mult_0_350  = SHARE((!Xd_0__inst_mult_0_528  & (Xd_0__inst_mult_0_532  & Xd_0__inst_mult_0_536 )) # (Xd_0__inst_mult_0_528  & ((Xd_0__inst_mult_0_536 ) # (Xd_0__inst_mult_0_532 ))))

	.dataa(!Xd_0__inst_mult_0_528 ),
	.datab(!Xd_0__inst_mult_0_532 ),
	.datac(!Xd_0__inst_mult_0_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_341 ),
	.sharein(Xd_0__inst_mult_0_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_348 ),
	.cout(Xd_0__inst_mult_0_349 ),
	.shareout(Xd_0__inst_mult_0_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_111 (
// Equation(s):
// Xd_0__inst_mult_1_344  = SUM(( !Xd_0__inst_mult_1_524  $ (((!din_b[16]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_338  ) + ( Xd_0__inst_mult_1_337  ))
// Xd_0__inst_mult_1_345  = CARRY(( !Xd_0__inst_mult_1_524  $ (((!din_b[16]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_338  ) + ( Xd_0__inst_mult_1_337  ))
// Xd_0__inst_mult_1_346  = SHARE((din_b[16] & (din_a[22] & Xd_0__inst_mult_1_524 )))

	.dataa(!din_b[16]),
	.datab(!din_a[22]),
	.datac(!Xd_0__inst_mult_1_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_337 ),
	.sharein(Xd_0__inst_mult_1_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_344 ),
	.cout(Xd_0__inst_mult_1_345 ),
	.shareout(Xd_0__inst_mult_1_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_112 (
// Equation(s):
// Xd_0__inst_mult_1_348  = SUM(( !Xd_0__inst_mult_1_528  $ (!Xd_0__inst_mult_1_532  $ (Xd_0__inst_mult_1_536 )) ) + ( Xd_0__inst_mult_1_342  ) + ( Xd_0__inst_mult_1_341  ))
// Xd_0__inst_mult_1_349  = CARRY(( !Xd_0__inst_mult_1_528  $ (!Xd_0__inst_mult_1_532  $ (Xd_0__inst_mult_1_536 )) ) + ( Xd_0__inst_mult_1_342  ) + ( Xd_0__inst_mult_1_341  ))
// Xd_0__inst_mult_1_350  = SHARE((!Xd_0__inst_mult_1_528  & (Xd_0__inst_mult_1_532  & Xd_0__inst_mult_1_536 )) # (Xd_0__inst_mult_1_528  & ((Xd_0__inst_mult_1_536 ) # (Xd_0__inst_mult_1_532 ))))

	.dataa(!Xd_0__inst_mult_1_528 ),
	.datab(!Xd_0__inst_mult_1_532 ),
	.datac(!Xd_0__inst_mult_1_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_341 ),
	.sharein(Xd_0__inst_mult_1_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_348 ),
	.cout(Xd_0__inst_mult_1_349 ),
	.shareout(Xd_0__inst_mult_1_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_12_118 (
// Equation(s):
// Xd_0__inst_mult_12_384  = SUM(( !Xd_0__inst_mult_12_556  $ (!Xd_0__inst_mult_12_272  $ (Xd_0__inst_mult_14_540 )) ) + ( Xd_0__inst_mult_12_382  ) + ( Xd_0__inst_mult_12_381  ))
// Xd_0__inst_mult_12_385  = CARRY(( !Xd_0__inst_mult_12_556  $ (!Xd_0__inst_mult_12_272  $ (Xd_0__inst_mult_14_540 )) ) + ( Xd_0__inst_mult_12_382  ) + ( Xd_0__inst_mult_12_381  ))
// Xd_0__inst_mult_12_386  = SHARE((!Xd_0__inst_mult_12_556  & (Xd_0__inst_mult_12_272  & Xd_0__inst_mult_14_540 )) # (Xd_0__inst_mult_12_556  & ((Xd_0__inst_mult_14_540 ) # (Xd_0__inst_mult_12_272 ))))

	.dataa(!Xd_0__inst_mult_12_556 ),
	.datab(!Xd_0__inst_mult_12_272 ),
	.datac(!Xd_0__inst_mult_14_540 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_381 ),
	.sharein(Xd_0__inst_mult_12_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_384 ),
	.cout(Xd_0__inst_mult_12_385 ),
	.shareout(Xd_0__inst_mult_12_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_13_116 (
// Equation(s):
// Xd_0__inst_mult_13_364  = SUM(( !Xd_0__inst_mult_13_540  $ (!Xd_0__inst_mult_13_544  $ (Xd_0__inst_mult_1_540 )) ) + ( Xd_0__inst_mult_13_362  ) + ( Xd_0__inst_mult_13_361  ))
// Xd_0__inst_mult_13_365  = CARRY(( !Xd_0__inst_mult_13_540  $ (!Xd_0__inst_mult_13_544  $ (Xd_0__inst_mult_1_540 )) ) + ( Xd_0__inst_mult_13_362  ) + ( Xd_0__inst_mult_13_361  ))
// Xd_0__inst_mult_13_366  = SHARE((!Xd_0__inst_mult_13_540  & (Xd_0__inst_mult_13_544  & Xd_0__inst_mult_1_540 )) # (Xd_0__inst_mult_13_540  & ((Xd_0__inst_mult_1_540 ) # (Xd_0__inst_mult_13_544 ))))

	.dataa(!Xd_0__inst_mult_13_540 ),
	.datab(!Xd_0__inst_mult_13_544 ),
	.datac(!Xd_0__inst_mult_1_540 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_361 ),
	.sharein(Xd_0__inst_mult_13_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_364 ),
	.cout(Xd_0__inst_mult_13_365 ),
	.shareout(Xd_0__inst_mult_13_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_14_120 (
// Equation(s):
// Xd_0__inst_mult_14_380  = SUM(( !Xd_0__inst_mult_14_544  $ (!Xd_0__inst_mult_14_548  $ (Xd_0__inst_mult_15_560 )) ) + ( Xd_0__inst_mult_14_378  ) + ( Xd_0__inst_mult_14_377  ))
// Xd_0__inst_mult_14_381  = CARRY(( !Xd_0__inst_mult_14_544  $ (!Xd_0__inst_mult_14_548  $ (Xd_0__inst_mult_15_560 )) ) + ( Xd_0__inst_mult_14_378  ) + ( Xd_0__inst_mult_14_377  ))
// Xd_0__inst_mult_14_382  = SHARE((!Xd_0__inst_mult_14_544  & (Xd_0__inst_mult_14_548  & Xd_0__inst_mult_15_560 )) # (Xd_0__inst_mult_14_544  & ((Xd_0__inst_mult_15_560 ) # (Xd_0__inst_mult_14_548 ))))

	.dataa(!Xd_0__inst_mult_14_544 ),
	.datab(!Xd_0__inst_mult_14_548 ),
	.datac(!Xd_0__inst_mult_15_560 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_377 ),
	.sharein(Xd_0__inst_mult_14_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_380 ),
	.cout(Xd_0__inst_mult_14_381 ),
	.shareout(Xd_0__inst_mult_14_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_15_122 (
// Equation(s):
// Xd_0__inst_mult_15_388  = SUM(( !Xd_0__inst_mult_15_564  $ (!Xd_0__inst_mult_15_268  $ (Xd_0__inst_mult_14_552 )) ) + ( Xd_0__inst_mult_15_386  ) + ( Xd_0__inst_mult_15_385  ))
// Xd_0__inst_mult_15_389  = CARRY(( !Xd_0__inst_mult_15_564  $ (!Xd_0__inst_mult_15_268  $ (Xd_0__inst_mult_14_552 )) ) + ( Xd_0__inst_mult_15_386  ) + ( Xd_0__inst_mult_15_385  ))
// Xd_0__inst_mult_15_390  = SHARE((!Xd_0__inst_mult_15_564  & (Xd_0__inst_mult_15_268  & Xd_0__inst_mult_14_552 )) # (Xd_0__inst_mult_15_564  & ((Xd_0__inst_mult_14_552 ) # (Xd_0__inst_mult_15_268 ))))

	.dataa(!Xd_0__inst_mult_15_564 ),
	.datab(!Xd_0__inst_mult_15_268 ),
	.datac(!Xd_0__inst_mult_14_552 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_385 ),
	.sharein(Xd_0__inst_mult_15_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_388 ),
	.cout(Xd_0__inst_mult_15_389 ),
	.shareout(Xd_0__inst_mult_15_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_10_112 (
// Equation(s):
// Xd_0__inst_mult_10_360  = SUM(( !Xd_0__inst_mult_10_536  $ (!Xd_0__inst_mult_10_540  $ (Xd_0__inst_mult_0_540 )) ) + ( Xd_0__inst_mult_10_358  ) + ( Xd_0__inst_mult_10_357  ))
// Xd_0__inst_mult_10_361  = CARRY(( !Xd_0__inst_mult_10_536  $ (!Xd_0__inst_mult_10_540  $ (Xd_0__inst_mult_0_540 )) ) + ( Xd_0__inst_mult_10_358  ) + ( Xd_0__inst_mult_10_357  ))
// Xd_0__inst_mult_10_362  = SHARE((!Xd_0__inst_mult_10_536  & (Xd_0__inst_mult_10_540  & Xd_0__inst_mult_0_540 )) # (Xd_0__inst_mult_10_536  & ((Xd_0__inst_mult_0_540 ) # (Xd_0__inst_mult_10_540 ))))

	.dataa(!Xd_0__inst_mult_10_536 ),
	.datab(!Xd_0__inst_mult_10_540 ),
	.datac(!Xd_0__inst_mult_0_540 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_357 ),
	.sharein(Xd_0__inst_mult_10_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_360 ),
	.cout(Xd_0__inst_mult_10_361 ),
	.shareout(Xd_0__inst_mult_10_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_11_116 (
// Equation(s):
// Xd_0__inst_mult_11_364  = SUM(( !Xd_0__inst_mult_11_540  $ (!Xd_0__inst_mult_11_544  $ (Xd_0__inst_mult_3_536 )) ) + ( Xd_0__inst_mult_11_362  ) + ( Xd_0__inst_mult_11_361  ))
// Xd_0__inst_mult_11_365  = CARRY(( !Xd_0__inst_mult_11_540  $ (!Xd_0__inst_mult_11_544  $ (Xd_0__inst_mult_3_536 )) ) + ( Xd_0__inst_mult_11_362  ) + ( Xd_0__inst_mult_11_361  ))
// Xd_0__inst_mult_11_366  = SHARE((!Xd_0__inst_mult_11_540  & (Xd_0__inst_mult_11_544  & Xd_0__inst_mult_3_536 )) # (Xd_0__inst_mult_11_540  & ((Xd_0__inst_mult_3_536 ) # (Xd_0__inst_mult_11_544 ))))

	.dataa(!Xd_0__inst_mult_11_540 ),
	.datab(!Xd_0__inst_mult_11_544 ),
	.datac(!Xd_0__inst_mult_3_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_361 ),
	.sharein(Xd_0__inst_mult_11_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_364 ),
	.cout(Xd_0__inst_mult_11_365 ),
	.shareout(Xd_0__inst_mult_11_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_8_116 (
// Equation(s):
// Xd_0__inst_mult_8_364  = SUM(( !Xd_0__inst_mult_8_540  $ (!Xd_0__inst_mult_8_544  $ (Xd_0__inst_mult_2_540 )) ) + ( Xd_0__inst_mult_8_362  ) + ( Xd_0__inst_mult_8_361  ))
// Xd_0__inst_mult_8_365  = CARRY(( !Xd_0__inst_mult_8_540  $ (!Xd_0__inst_mult_8_544  $ (Xd_0__inst_mult_2_540 )) ) + ( Xd_0__inst_mult_8_362  ) + ( Xd_0__inst_mult_8_361  ))
// Xd_0__inst_mult_8_366  = SHARE((!Xd_0__inst_mult_8_540  & (Xd_0__inst_mult_8_544  & Xd_0__inst_mult_2_540 )) # (Xd_0__inst_mult_8_540  & ((Xd_0__inst_mult_2_540 ) # (Xd_0__inst_mult_8_544 ))))

	.dataa(!Xd_0__inst_mult_8_540 ),
	.datab(!Xd_0__inst_mult_8_544 ),
	.datac(!Xd_0__inst_mult_2_540 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_361 ),
	.sharein(Xd_0__inst_mult_8_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_364 ),
	.cout(Xd_0__inst_mult_8_365 ),
	.shareout(Xd_0__inst_mult_8_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_9_112 (
// Equation(s):
// Xd_0__inst_mult_9_360  = SUM(( !Xd_0__inst_mult_9_536  $ (!Xd_0__inst_mult_9_540  $ (Xd_0__inst_mult_1_544 )) ) + ( Xd_0__inst_mult_9_358  ) + ( Xd_0__inst_mult_9_357  ))
// Xd_0__inst_mult_9_361  = CARRY(( !Xd_0__inst_mult_9_536  $ (!Xd_0__inst_mult_9_540  $ (Xd_0__inst_mult_1_544 )) ) + ( Xd_0__inst_mult_9_358  ) + ( Xd_0__inst_mult_9_357  ))
// Xd_0__inst_mult_9_362  = SHARE((!Xd_0__inst_mult_9_536  & (Xd_0__inst_mult_9_540  & Xd_0__inst_mult_1_544 )) # (Xd_0__inst_mult_9_536  & ((Xd_0__inst_mult_1_544 ) # (Xd_0__inst_mult_9_540 ))))

	.dataa(!Xd_0__inst_mult_9_536 ),
	.datab(!Xd_0__inst_mult_9_540 ),
	.datac(!Xd_0__inst_mult_1_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_357 ),
	.sharein(Xd_0__inst_mult_9_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_360 ),
	.cout(Xd_0__inst_mult_9_361 ),
	.shareout(Xd_0__inst_mult_9_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_112 (
// Equation(s):
// Xd_0__inst_mult_6_360  = SUM(( !Xd_0__inst_mult_6_536  $ (!Xd_0__inst_mult_6_540  $ (Xd_0__inst_mult_5_536 )) ) + ( Xd_0__inst_mult_6_358  ) + ( Xd_0__inst_mult_6_357  ))
// Xd_0__inst_mult_6_361  = CARRY(( !Xd_0__inst_mult_6_536  $ (!Xd_0__inst_mult_6_540  $ (Xd_0__inst_mult_5_536 )) ) + ( Xd_0__inst_mult_6_358  ) + ( Xd_0__inst_mult_6_357  ))
// Xd_0__inst_mult_6_362  = SHARE((!Xd_0__inst_mult_6_536  & (Xd_0__inst_mult_6_540  & Xd_0__inst_mult_5_536 )) # (Xd_0__inst_mult_6_536  & ((Xd_0__inst_mult_5_536 ) # (Xd_0__inst_mult_6_540 ))))

	.dataa(!Xd_0__inst_mult_6_536 ),
	.datab(!Xd_0__inst_mult_6_540 ),
	.datac(!Xd_0__inst_mult_5_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_357 ),
	.sharein(Xd_0__inst_mult_6_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_360 ),
	.cout(Xd_0__inst_mult_6_361 ),
	.shareout(Xd_0__inst_mult_6_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_109 (
// Equation(s):
// Xd_0__inst_mult_7_348  = SUM(( GND ) + ( Xd_0__inst_mult_7_342  ) + ( Xd_0__inst_mult_7_341  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_341 ),
	.sharein(Xd_0__inst_mult_7_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_348 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_110 (
// Equation(s):
// Xd_0__inst_mult_7_352  = SUM(( !Xd_0__inst_mult_7_536  $ (!Xd_0__inst_mult_7_540  $ (Xd_0__inst_mult_7_544 )) ) + ( Xd_0__inst_mult_7_346  ) + ( Xd_0__inst_mult_7_345  ))
// Xd_0__inst_mult_7_353  = CARRY(( !Xd_0__inst_mult_7_536  $ (!Xd_0__inst_mult_7_540  $ (Xd_0__inst_mult_7_544 )) ) + ( Xd_0__inst_mult_7_346  ) + ( Xd_0__inst_mult_7_345  ))
// Xd_0__inst_mult_7_354  = SHARE((!Xd_0__inst_mult_7_536  & (Xd_0__inst_mult_7_540  & Xd_0__inst_mult_7_544 )) # (Xd_0__inst_mult_7_536  & ((Xd_0__inst_mult_7_544 ) # (Xd_0__inst_mult_7_540 ))))

	.dataa(!Xd_0__inst_mult_7_536 ),
	.datab(!Xd_0__inst_mult_7_540 ),
	.datac(!Xd_0__inst_mult_7_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_345 ),
	.sharein(Xd_0__inst_mult_7_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_352 ),
	.cout(Xd_0__inst_mult_7_353 ),
	.shareout(Xd_0__inst_mult_7_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_121 (
// Equation(s):
// Xd_0__inst_mult_4_384  = SUM(( GND ) + ( Xd_0__inst_mult_4_378  ) + ( Xd_0__inst_mult_4_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_377 ),
	.sharein(Xd_0__inst_mult_4_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_384 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_122 (
// Equation(s):
// Xd_0__inst_mult_4_388  = SUM(( !Xd_0__inst_mult_4_560  $ (!Xd_0__inst_mult_4_188  $ (Xd_0__inst_mult_6_544 )) ) + ( Xd_0__inst_mult_4_382  ) + ( Xd_0__inst_mult_4_381  ))
// Xd_0__inst_mult_4_389  = CARRY(( !Xd_0__inst_mult_4_560  $ (!Xd_0__inst_mult_4_188  $ (Xd_0__inst_mult_6_544 )) ) + ( Xd_0__inst_mult_4_382  ) + ( Xd_0__inst_mult_4_381  ))
// Xd_0__inst_mult_4_390  = SHARE((!Xd_0__inst_mult_4_560  & (Xd_0__inst_mult_4_188  & Xd_0__inst_mult_6_544 )) # (Xd_0__inst_mult_4_560  & ((Xd_0__inst_mult_6_544 ) # (Xd_0__inst_mult_4_188 ))))

	.dataa(!Xd_0__inst_mult_4_560 ),
	.datab(!Xd_0__inst_mult_4_188 ),
	.datac(!Xd_0__inst_mult_6_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_381 ),
	.sharein(Xd_0__inst_mult_4_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_388 ),
	.cout(Xd_0__inst_mult_4_389 ),
	.shareout(Xd_0__inst_mult_4_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_109 (
// Equation(s):
// Xd_0__inst_mult_5_348  = SUM(( GND ) + ( Xd_0__inst_mult_5_342  ) + ( Xd_0__inst_mult_5_341  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_341 ),
	.sharein(Xd_0__inst_mult_5_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_348 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_110 (
// Equation(s):
// Xd_0__inst_mult_5_352  = SUM(( !Xd_0__inst_mult_5_540  $ (!Xd_0__inst_mult_5_544  $ (Xd_0__inst_mult_9_544 )) ) + ( Xd_0__inst_mult_5_346  ) + ( Xd_0__inst_mult_5_345  ))
// Xd_0__inst_mult_5_353  = CARRY(( !Xd_0__inst_mult_5_540  $ (!Xd_0__inst_mult_5_544  $ (Xd_0__inst_mult_9_544 )) ) + ( Xd_0__inst_mult_5_346  ) + ( Xd_0__inst_mult_5_345  ))
// Xd_0__inst_mult_5_354  = SHARE((!Xd_0__inst_mult_5_540  & (Xd_0__inst_mult_5_544  & Xd_0__inst_mult_9_544 )) # (Xd_0__inst_mult_5_540  & ((Xd_0__inst_mult_9_544 ) # (Xd_0__inst_mult_5_544 ))))

	.dataa(!Xd_0__inst_mult_5_540 ),
	.datab(!Xd_0__inst_mult_5_544 ),
	.datac(!Xd_0__inst_mult_9_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_345 ),
	.sharein(Xd_0__inst_mult_5_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_352 ),
	.cout(Xd_0__inst_mult_5_353 ),
	.shareout(Xd_0__inst_mult_5_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_113 (
// Equation(s):
// Xd_0__inst_mult_2_352  = SUM(( GND ) + ( Xd_0__inst_mult_2_346  ) + ( Xd_0__inst_mult_2_345  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_345 ),
	.sharein(Xd_0__inst_mult_2_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_352 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_114 (
// Equation(s):
// Xd_0__inst_mult_2_356  = SUM(( !Xd_0__inst_mult_2_544  $ (!Xd_0__inst_mult_2_548  $ (Xd_0__inst_mult_13_548 )) ) + ( Xd_0__inst_mult_2_350  ) + ( Xd_0__inst_mult_2_349  ))
// Xd_0__inst_mult_2_357  = CARRY(( !Xd_0__inst_mult_2_544  $ (!Xd_0__inst_mult_2_548  $ (Xd_0__inst_mult_13_548 )) ) + ( Xd_0__inst_mult_2_350  ) + ( Xd_0__inst_mult_2_349  ))
// Xd_0__inst_mult_2_358  = SHARE((!Xd_0__inst_mult_2_544  & (Xd_0__inst_mult_2_548  & Xd_0__inst_mult_13_548 )) # (Xd_0__inst_mult_2_544  & ((Xd_0__inst_mult_13_548 ) # (Xd_0__inst_mult_2_548 ))))

	.dataa(!Xd_0__inst_mult_2_544 ),
	.datab(!Xd_0__inst_mult_2_548 ),
	.datac(!Xd_0__inst_mult_13_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_349 ),
	.sharein(Xd_0__inst_mult_2_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_356 ),
	.cout(Xd_0__inst_mult_2_357 ),
	.shareout(Xd_0__inst_mult_2_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_109 (
// Equation(s):
// Xd_0__inst_mult_3_348  = SUM(( GND ) + ( Xd_0__inst_mult_3_342  ) + ( Xd_0__inst_mult_3_341  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_341 ),
	.sharein(Xd_0__inst_mult_3_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_348 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_110 (
// Equation(s):
// Xd_0__inst_mult_3_352  = SUM(( !Xd_0__inst_mult_3_540  $ (!Xd_0__inst_mult_3_544  $ (Xd_0__inst_mult_8_548 )) ) + ( Xd_0__inst_mult_3_346  ) + ( Xd_0__inst_mult_3_345  ))
// Xd_0__inst_mult_3_353  = CARRY(( !Xd_0__inst_mult_3_540  $ (!Xd_0__inst_mult_3_544  $ (Xd_0__inst_mult_8_548 )) ) + ( Xd_0__inst_mult_3_346  ) + ( Xd_0__inst_mult_3_345  ))
// Xd_0__inst_mult_3_354  = SHARE((!Xd_0__inst_mult_3_540  & (Xd_0__inst_mult_3_544  & Xd_0__inst_mult_8_548 )) # (Xd_0__inst_mult_3_540  & ((Xd_0__inst_mult_8_548 ) # (Xd_0__inst_mult_3_544 ))))

	.dataa(!Xd_0__inst_mult_3_540 ),
	.datab(!Xd_0__inst_mult_3_544 ),
	.datac(!Xd_0__inst_mult_8_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_345 ),
	.sharein(Xd_0__inst_mult_3_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_352 ),
	.cout(Xd_0__inst_mult_3_353 ),
	.shareout(Xd_0__inst_mult_3_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_113 (
// Equation(s):
// Xd_0__inst_mult_0_352  = SUM(( GND ) + ( Xd_0__inst_mult_0_346  ) + ( Xd_0__inst_mult_0_345  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_345 ),
	.sharein(Xd_0__inst_mult_0_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_352 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_114 (
// Equation(s):
// Xd_0__inst_mult_0_356  = SUM(( !Xd_0__inst_mult_0_544  $ (!Xd_0__inst_mult_0_548  $ (Xd_0__inst_mult_11_548 )) ) + ( Xd_0__inst_mult_0_350  ) + ( Xd_0__inst_mult_0_349  ))
// Xd_0__inst_mult_0_357  = CARRY(( !Xd_0__inst_mult_0_544  $ (!Xd_0__inst_mult_0_548  $ (Xd_0__inst_mult_11_548 )) ) + ( Xd_0__inst_mult_0_350  ) + ( Xd_0__inst_mult_0_349  ))
// Xd_0__inst_mult_0_358  = SHARE((!Xd_0__inst_mult_0_544  & (Xd_0__inst_mult_0_548  & Xd_0__inst_mult_11_548 )) # (Xd_0__inst_mult_0_544  & ((Xd_0__inst_mult_11_548 ) # (Xd_0__inst_mult_0_548 ))))

	.dataa(!Xd_0__inst_mult_0_544 ),
	.datab(!Xd_0__inst_mult_0_548 ),
	.datac(!Xd_0__inst_mult_11_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_349 ),
	.sharein(Xd_0__inst_mult_0_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_356 ),
	.cout(Xd_0__inst_mult_0_357 ),
	.shareout(Xd_0__inst_mult_0_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_113 (
// Equation(s):
// Xd_0__inst_mult_1_352  = SUM(( GND ) + ( Xd_0__inst_mult_1_346  ) + ( Xd_0__inst_mult_1_345  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_345 ),
	.sharein(Xd_0__inst_mult_1_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_352 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_114 (
// Equation(s):
// Xd_0__inst_mult_1_356  = SUM(( !Xd_0__inst_mult_1_548  $ (!Xd_0__inst_mult_1_552  $ (Xd_0__inst_mult_10_544 )) ) + ( Xd_0__inst_mult_1_350  ) + ( Xd_0__inst_mult_1_349  ))
// Xd_0__inst_mult_1_357  = CARRY(( !Xd_0__inst_mult_1_548  $ (!Xd_0__inst_mult_1_552  $ (Xd_0__inst_mult_10_544 )) ) + ( Xd_0__inst_mult_1_350  ) + ( Xd_0__inst_mult_1_349  ))
// Xd_0__inst_mult_1_358  = SHARE((!Xd_0__inst_mult_1_548  & (Xd_0__inst_mult_1_552  & Xd_0__inst_mult_10_544 )) # (Xd_0__inst_mult_1_548  & ((Xd_0__inst_mult_10_544 ) # (Xd_0__inst_mult_1_552 ))))

	.dataa(!Xd_0__inst_mult_1_548 ),
	.datab(!Xd_0__inst_mult_1_552 ),
	.datac(!Xd_0__inst_mult_10_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_349 ),
	.sharein(Xd_0__inst_mult_1_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_356 ),
	.cout(Xd_0__inst_mult_1_357 ),
	.shareout(Xd_0__inst_mult_1_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_119 (
// Equation(s):
// Xd_0__inst_mult_12_388  = SUM(( !Xd_0__inst_mult_12_560  $ (!Xd_0__inst_mult_12_188 ) ) + ( Xd_0__inst_mult_12_386  ) + ( Xd_0__inst_mult_12_385  ))
// Xd_0__inst_mult_12_389  = CARRY(( !Xd_0__inst_mult_12_560  $ (!Xd_0__inst_mult_12_188 ) ) + ( Xd_0__inst_mult_12_386  ) + ( Xd_0__inst_mult_12_385  ))
// Xd_0__inst_mult_12_390  = SHARE((Xd_0__inst_mult_12_560  & Xd_0__inst_mult_12_188 ))

	.dataa(!Xd_0__inst_mult_12_560 ),
	.datab(!Xd_0__inst_mult_12_188 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_385 ),
	.sharein(Xd_0__inst_mult_12_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_388 ),
	.cout(Xd_0__inst_mult_12_389 ),
	.shareout(Xd_0__inst_mult_12_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_47 (
// Equation(s):
// Xd_0__inst_mult_12_47_sumout  = SUM(( (din_a[154] & din_b[150]) ) + ( Xd_0__inst_mult_11_53  ) + ( Xd_0__inst_mult_11_52  ))
// Xd_0__inst_mult_12_48  = CARRY(( (din_a[154] & din_b[150]) ) + ( Xd_0__inst_mult_11_53  ) + ( Xd_0__inst_mult_11_52  ))
// Xd_0__inst_mult_12_49  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[150]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_52 ),
	.sharein(Xd_0__inst_mult_11_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_47_sumout ),
	.cout(Xd_0__inst_mult_12_48 ),
	.shareout(Xd_0__inst_mult_12_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_117 (
// Equation(s):
// Xd_0__inst_mult_13_368  = SUM(( !Xd_0__inst_mult_13_552  $ (!Xd_0__inst_mult_13_556 ) ) + ( Xd_0__inst_mult_13_366  ) + ( Xd_0__inst_mult_13_365  ))
// Xd_0__inst_mult_13_369  = CARRY(( !Xd_0__inst_mult_13_552  $ (!Xd_0__inst_mult_13_556 ) ) + ( Xd_0__inst_mult_13_366  ) + ( Xd_0__inst_mult_13_365  ))
// Xd_0__inst_mult_13_370  = SHARE((Xd_0__inst_mult_13_552  & Xd_0__inst_mult_13_556 ))

	.dataa(!Xd_0__inst_mult_13_552 ),
	.datab(!Xd_0__inst_mult_13_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_365 ),
	.sharein(Xd_0__inst_mult_13_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_368 ),
	.cout(Xd_0__inst_mult_13_369 ),
	.shareout(Xd_0__inst_mult_13_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_43 (
// Equation(s):
// Xd_0__inst_mult_13_43_sumout  = SUM(( (din_a[166] & din_b[162]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_44  = CARRY(( (din_a[166] & din_b[162]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_45  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[162]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_13_43_sumout ),
	.cout(Xd_0__inst_mult_13_44 ),
	.shareout(Xd_0__inst_mult_13_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_121 (
// Equation(s):
// Xd_0__inst_mult_14_384  = SUM(( !Xd_0__inst_mult_14_556  $ (!Xd_0__inst_mult_14_560 ) ) + ( Xd_0__inst_mult_14_382  ) + ( Xd_0__inst_mult_14_381  ))
// Xd_0__inst_mult_14_385  = CARRY(( !Xd_0__inst_mult_14_556  $ (!Xd_0__inst_mult_14_560 ) ) + ( Xd_0__inst_mult_14_382  ) + ( Xd_0__inst_mult_14_381  ))
// Xd_0__inst_mult_14_386  = SHARE((Xd_0__inst_mult_14_556  & Xd_0__inst_mult_14_560 ))

	.dataa(!Xd_0__inst_mult_14_556 ),
	.datab(!Xd_0__inst_mult_14_560 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_381 ),
	.sharein(Xd_0__inst_mult_14_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_384 ),
	.cout(Xd_0__inst_mult_14_385 ),
	.shareout(Xd_0__inst_mult_14_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_123 (
// Equation(s):
// Xd_0__inst_mult_15_392  = SUM(( !Xd_0__inst_mult_15_568  $ (!Xd_0__inst_mult_15_188 ) ) + ( Xd_0__inst_mult_15_390  ) + ( Xd_0__inst_mult_15_389  ))
// Xd_0__inst_mult_15_393  = CARRY(( !Xd_0__inst_mult_15_568  $ (!Xd_0__inst_mult_15_188 ) ) + ( Xd_0__inst_mult_15_390  ) + ( Xd_0__inst_mult_15_389  ))
// Xd_0__inst_mult_15_394  = SHARE((Xd_0__inst_mult_15_568  & Xd_0__inst_mult_15_188 ))

	.dataa(!Xd_0__inst_mult_15_568 ),
	.datab(!Xd_0__inst_mult_15_188 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_389 ),
	.sharein(Xd_0__inst_mult_15_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_392 ),
	.cout(Xd_0__inst_mult_15_393 ),
	.shareout(Xd_0__inst_mult_15_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_47 (
// Equation(s):
// Xd_0__inst_mult_15_47_sumout  = SUM(( (din_a[190] & din_b[186]) ) + ( Xd_0__inst_mult_12_49  ) + ( Xd_0__inst_mult_12_48  ))
// Xd_0__inst_mult_15_48  = CARRY(( (din_a[190] & din_b[186]) ) + ( Xd_0__inst_mult_12_49  ) + ( Xd_0__inst_mult_12_48  ))
// Xd_0__inst_mult_15_49  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[186]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_48 ),
	.sharein(Xd_0__inst_mult_12_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_47_sumout ),
	.cout(Xd_0__inst_mult_15_48 ),
	.shareout(Xd_0__inst_mult_15_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_113 (
// Equation(s):
// Xd_0__inst_mult_10_364  = SUM(( !Xd_0__inst_mult_10_548  $ (!Xd_0__inst_mult_10_552 ) ) + ( Xd_0__inst_mult_10_362  ) + ( Xd_0__inst_mult_10_361  ))
// Xd_0__inst_mult_10_365  = CARRY(( !Xd_0__inst_mult_10_548  $ (!Xd_0__inst_mult_10_552 ) ) + ( Xd_0__inst_mult_10_362  ) + ( Xd_0__inst_mult_10_361  ))
// Xd_0__inst_mult_10_366  = SHARE((Xd_0__inst_mult_10_548  & Xd_0__inst_mult_10_552 ))

	.dataa(!Xd_0__inst_mult_10_548 ),
	.datab(!Xd_0__inst_mult_10_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_361 ),
	.sharein(Xd_0__inst_mult_10_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_364 ),
	.cout(Xd_0__inst_mult_10_365 ),
	.shareout(Xd_0__inst_mult_10_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_115 (
// Equation(s):
// Xd_0__inst_mult_0_360  = SUM(( (din_a[130] & din_b[126]) ) + ( Xd_0__inst_mult_11_41  ) + ( Xd_0__inst_mult_11_40  ))
// Xd_0__inst_mult_0_361  = CARRY(( (din_a[130] & din_b[126]) ) + ( Xd_0__inst_mult_11_41  ) + ( Xd_0__inst_mult_11_40  ))
// Xd_0__inst_mult_0_362  = SHARE(Xd_0__inst_mult_0_384 )

	.dataa(!din_a[130]),
	.datab(!din_b[126]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_0_384 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_40 ),
	.sharein(Xd_0__inst_mult_11_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_360 ),
	.cout(Xd_0__inst_mult_0_361 ),
	.shareout(Xd_0__inst_mult_0_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_117 (
// Equation(s):
// Xd_0__inst_mult_11_368  = SUM(( !Xd_0__inst_mult_11_552  $ (!Xd_0__inst_mult_11_556 ) ) + ( Xd_0__inst_mult_11_366  ) + ( Xd_0__inst_mult_11_365  ))
// Xd_0__inst_mult_11_369  = CARRY(( !Xd_0__inst_mult_11_552  $ (!Xd_0__inst_mult_11_556 ) ) + ( Xd_0__inst_mult_11_366  ) + ( Xd_0__inst_mult_11_365  ))
// Xd_0__inst_mult_11_370  = SHARE((Xd_0__inst_mult_11_552  & Xd_0__inst_mult_11_556 ))

	.dataa(!Xd_0__inst_mult_11_552 ),
	.datab(!Xd_0__inst_mult_11_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_365 ),
	.sharein(Xd_0__inst_mult_11_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_368 ),
	.cout(Xd_0__inst_mult_11_369 ),
	.shareout(Xd_0__inst_mult_11_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_39 (
// Equation(s):
// Xd_0__inst_mult_11_39_sumout  = SUM(( (din_a[142] & din_b[138]) ) + ( Xd_0__inst_mult_8_49  ) + ( Xd_0__inst_mult_8_48  ))
// Xd_0__inst_mult_11_40  = CARRY(( (din_a[142] & din_b[138]) ) + ( Xd_0__inst_mult_8_49  ) + ( Xd_0__inst_mult_8_48  ))
// Xd_0__inst_mult_11_41  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[138]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_48 ),
	.sharein(Xd_0__inst_mult_8_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_39_sumout ),
	.cout(Xd_0__inst_mult_11_40 ),
	.shareout(Xd_0__inst_mult_11_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_117 (
// Equation(s):
// Xd_0__inst_mult_8_368  = SUM(( !Xd_0__inst_mult_8_552  $ (!Xd_0__inst_mult_8_556 ) ) + ( Xd_0__inst_mult_8_366  ) + ( Xd_0__inst_mult_8_365  ))
// Xd_0__inst_mult_8_369  = CARRY(( !Xd_0__inst_mult_8_552  $ (!Xd_0__inst_mult_8_556 ) ) + ( Xd_0__inst_mult_8_366  ) + ( Xd_0__inst_mult_8_365  ))
// Xd_0__inst_mult_8_370  = SHARE((Xd_0__inst_mult_8_552  & Xd_0__inst_mult_8_556 ))

	.dataa(!Xd_0__inst_mult_8_552 ),
	.datab(!Xd_0__inst_mult_8_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_365 ),
	.sharein(Xd_0__inst_mult_8_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_368 ),
	.cout(Xd_0__inst_mult_8_369 ),
	.shareout(Xd_0__inst_mult_8_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_47 (
// Equation(s):
// Xd_0__inst_mult_8_47_sumout  = SUM(( (din_a[106] & din_b[102]) ) + ( Xd_0__inst_mult_9_41  ) + ( Xd_0__inst_mult_9_40  ))
// Xd_0__inst_mult_8_48  = CARRY(( (din_a[106] & din_b[102]) ) + ( Xd_0__inst_mult_9_41  ) + ( Xd_0__inst_mult_9_40  ))
// Xd_0__inst_mult_8_49  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[102]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_40 ),
	.sharein(Xd_0__inst_mult_9_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_47_sumout ),
	.cout(Xd_0__inst_mult_8_48 ),
	.shareout(Xd_0__inst_mult_8_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_113 (
// Equation(s):
// Xd_0__inst_mult_9_364  = SUM(( !Xd_0__inst_mult_9_548  $ (!Xd_0__inst_mult_9_552 ) ) + ( Xd_0__inst_mult_9_362  ) + ( Xd_0__inst_mult_9_361  ))
// Xd_0__inst_mult_9_365  = CARRY(( !Xd_0__inst_mult_9_548  $ (!Xd_0__inst_mult_9_552 ) ) + ( Xd_0__inst_mult_9_362  ) + ( Xd_0__inst_mult_9_361  ))
// Xd_0__inst_mult_9_366  = SHARE((Xd_0__inst_mult_9_548  & Xd_0__inst_mult_9_552 ))

	.dataa(!Xd_0__inst_mult_9_548 ),
	.datab(!Xd_0__inst_mult_9_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_361 ),
	.sharein(Xd_0__inst_mult_9_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_364 ),
	.cout(Xd_0__inst_mult_9_365 ),
	.shareout(Xd_0__inst_mult_9_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_39 (
// Equation(s):
// Xd_0__inst_mult_9_39_sumout  = SUM(( (din_a[118] & din_b[114]) ) + ( Xd_0__inst_mult_6_45  ) + ( Xd_0__inst_mult_6_44  ))
// Xd_0__inst_mult_9_40  = CARRY(( (din_a[118] & din_b[114]) ) + ( Xd_0__inst_mult_6_45  ) + ( Xd_0__inst_mult_6_44  ))
// Xd_0__inst_mult_9_41  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[114]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_44 ),
	.sharein(Xd_0__inst_mult_6_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_39_sumout ),
	.cout(Xd_0__inst_mult_9_40 ),
	.shareout(Xd_0__inst_mult_9_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_113 (
// Equation(s):
// Xd_0__inst_mult_6_364  = SUM(( !Xd_0__inst_mult_6_548  $ (!Xd_0__inst_mult_6_552 ) ) + ( Xd_0__inst_mult_6_362  ) + ( Xd_0__inst_mult_6_361  ))
// Xd_0__inst_mult_6_365  = CARRY(( !Xd_0__inst_mult_6_548  $ (!Xd_0__inst_mult_6_552 ) ) + ( Xd_0__inst_mult_6_362  ) + ( Xd_0__inst_mult_6_361  ))
// Xd_0__inst_mult_6_366  = SHARE((Xd_0__inst_mult_6_548  & Xd_0__inst_mult_6_552 ))

	.dataa(!Xd_0__inst_mult_6_548 ),
	.datab(!Xd_0__inst_mult_6_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_361 ),
	.sharein(Xd_0__inst_mult_6_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_364 ),
	.cout(Xd_0__inst_mult_6_365 ),
	.shareout(Xd_0__inst_mult_6_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_43 (
// Equation(s):
// Xd_0__inst_mult_6_43_sumout  = SUM(( (din_a[82] & din_b[78]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_44  = CARRY(( (din_a[82] & din_b[78]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_45  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[78]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_43_sumout ),
	.cout(Xd_0__inst_mult_6_44 ),
	.shareout(Xd_0__inst_mult_6_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_111 (
// Equation(s):
// Xd_0__inst_mult_7_356  = SUM(( !Xd_0__inst_mult_7_548  $ (!Xd_0__inst_mult_7_552 ) ) + ( Xd_0__inst_mult_7_354  ) + ( Xd_0__inst_mult_7_353  ))
// Xd_0__inst_mult_7_357  = CARRY(( !Xd_0__inst_mult_7_548  $ (!Xd_0__inst_mult_7_552 ) ) + ( Xd_0__inst_mult_7_354  ) + ( Xd_0__inst_mult_7_353  ))
// Xd_0__inst_mult_7_358  = SHARE((Xd_0__inst_mult_7_548  & Xd_0__inst_mult_7_552 ))

	.dataa(!Xd_0__inst_mult_7_548 ),
	.datab(!Xd_0__inst_mult_7_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_353 ),
	.sharein(Xd_0__inst_mult_7_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_356 ),
	.cout(Xd_0__inst_mult_7_357 ),
	.shareout(Xd_0__inst_mult_7_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_115 (
// Equation(s):
// Xd_0__inst_mult_1_360  = SUM(( (din_a[94] & din_b[90]) ) + ( Xd_0__inst_mult_4_41  ) + ( Xd_0__inst_mult_4_40  ))
// Xd_0__inst_mult_1_361  = CARRY(( (din_a[94] & din_b[90]) ) + ( Xd_0__inst_mult_4_41  ) + ( Xd_0__inst_mult_4_40  ))
// Xd_0__inst_mult_1_362  = SHARE(Xd_0__inst_mult_1_384 )

	.dataa(!din_a[94]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_1_384 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_40 ),
	.sharein(Xd_0__inst_mult_4_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_360 ),
	.cout(Xd_0__inst_mult_1_361 ),
	.shareout(Xd_0__inst_mult_1_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_123 (
// Equation(s):
// Xd_0__inst_mult_4_392  = SUM(( !Xd_0__inst_mult_4_564  $ (!Xd_0__inst_mult_4_184 ) ) + ( Xd_0__inst_mult_4_390  ) + ( Xd_0__inst_mult_4_389  ))
// Xd_0__inst_mult_4_393  = CARRY(( !Xd_0__inst_mult_4_564  $ (!Xd_0__inst_mult_4_184 ) ) + ( Xd_0__inst_mult_4_390  ) + ( Xd_0__inst_mult_4_389  ))
// Xd_0__inst_mult_4_394  = SHARE((Xd_0__inst_mult_4_564  & Xd_0__inst_mult_4_184 ))

	.dataa(!Xd_0__inst_mult_4_564 ),
	.datab(!Xd_0__inst_mult_4_184 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_389 ),
	.sharein(Xd_0__inst_mult_4_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_392 ),
	.cout(Xd_0__inst_mult_4_393 ),
	.shareout(Xd_0__inst_mult_4_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_39 (
// Equation(s):
// Xd_0__inst_mult_4_39_sumout  = SUM(( (din_a[58] & din_b[54]) ) + ( Xd_0__inst_mult_5_45  ) + ( Xd_0__inst_mult_5_44  ))
// Xd_0__inst_mult_4_40  = CARRY(( (din_a[58] & din_b[54]) ) + ( Xd_0__inst_mult_5_45  ) + ( Xd_0__inst_mult_5_44  ))
// Xd_0__inst_mult_4_41  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_44 ),
	.sharein(Xd_0__inst_mult_5_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_39_sumout ),
	.cout(Xd_0__inst_mult_4_40 ),
	.shareout(Xd_0__inst_mult_4_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_111 (
// Equation(s):
// Xd_0__inst_mult_5_356  = SUM(( !Xd_0__inst_mult_5_548  $ (!Xd_0__inst_mult_5_552 ) ) + ( Xd_0__inst_mult_5_354  ) + ( Xd_0__inst_mult_5_353  ))
// Xd_0__inst_mult_5_357  = CARRY(( !Xd_0__inst_mult_5_548  $ (!Xd_0__inst_mult_5_552 ) ) + ( Xd_0__inst_mult_5_354  ) + ( Xd_0__inst_mult_5_353  ))
// Xd_0__inst_mult_5_358  = SHARE((Xd_0__inst_mult_5_548  & Xd_0__inst_mult_5_552 ))

	.dataa(!Xd_0__inst_mult_5_548 ),
	.datab(!Xd_0__inst_mult_5_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_353 ),
	.sharein(Xd_0__inst_mult_5_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_356 ),
	.cout(Xd_0__inst_mult_5_357 ),
	.shareout(Xd_0__inst_mult_5_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_43 (
// Equation(s):
// Xd_0__inst_mult_5_43_sumout  = SUM(( (din_a[70] & din_b[66]) ) + ( Xd_0__inst_mult_2_45  ) + ( Xd_0__inst_mult_2_44  ))
// Xd_0__inst_mult_5_44  = CARRY(( (din_a[70] & din_b[66]) ) + ( Xd_0__inst_mult_2_45  ) + ( Xd_0__inst_mult_2_44  ))
// Xd_0__inst_mult_5_45  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[66]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_44 ),
	.sharein(Xd_0__inst_mult_2_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_43_sumout ),
	.cout(Xd_0__inst_mult_5_44 ),
	.shareout(Xd_0__inst_mult_5_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_115 (
// Equation(s):
// Xd_0__inst_mult_2_360  = SUM(( !Xd_0__inst_mult_2_552  $ (!Xd_0__inst_mult_2_556 ) ) + ( Xd_0__inst_mult_2_358  ) + ( Xd_0__inst_mult_2_357  ))
// Xd_0__inst_mult_2_361  = CARRY(( !Xd_0__inst_mult_2_552  $ (!Xd_0__inst_mult_2_556 ) ) + ( Xd_0__inst_mult_2_358  ) + ( Xd_0__inst_mult_2_357  ))
// Xd_0__inst_mult_2_362  = SHARE((Xd_0__inst_mult_2_552  & Xd_0__inst_mult_2_556 ))

	.dataa(!Xd_0__inst_mult_2_552 ),
	.datab(!Xd_0__inst_mult_2_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_357 ),
	.sharein(Xd_0__inst_mult_2_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_360 ),
	.cout(Xd_0__inst_mult_2_361 ),
	.shareout(Xd_0__inst_mult_2_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_43 (
// Equation(s):
// Xd_0__inst_mult_2_43_sumout  = SUM(( (din_a[34] & din_b[30]) ) + ( Xd_0__inst_mult_13_45  ) + ( Xd_0__inst_mult_13_44  ))
// Xd_0__inst_mult_2_44  = CARRY(( (din_a[34] & din_b[30]) ) + ( Xd_0__inst_mult_13_45  ) + ( Xd_0__inst_mult_13_44  ))
// Xd_0__inst_mult_2_45  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_44 ),
	.sharein(Xd_0__inst_mult_13_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_43_sumout ),
	.cout(Xd_0__inst_mult_2_44 ),
	.shareout(Xd_0__inst_mult_2_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_111 (
// Equation(s):
// Xd_0__inst_mult_3_356  = SUM(( !Xd_0__inst_mult_3_548  $ (!Xd_0__inst_mult_3_552 ) ) + ( Xd_0__inst_mult_3_354  ) + ( Xd_0__inst_mult_3_353  ))
// Xd_0__inst_mult_3_357  = CARRY(( !Xd_0__inst_mult_3_548  $ (!Xd_0__inst_mult_3_552 ) ) + ( Xd_0__inst_mult_3_354  ) + ( Xd_0__inst_mult_3_353  ))
// Xd_0__inst_mult_3_358  = SHARE((Xd_0__inst_mult_3_548  & Xd_0__inst_mult_3_552 ))

	.dataa(!Xd_0__inst_mult_3_548 ),
	.datab(!Xd_0__inst_mult_3_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_353 ),
	.sharein(Xd_0__inst_mult_3_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_356 ),
	.cout(Xd_0__inst_mult_3_357 ),
	.shareout(Xd_0__inst_mult_3_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_47 (
// Equation(s):
// Xd_0__inst_mult_3_47_sumout  = SUM(( (din_a[46] & din_b[42]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_48  = CARRY(( (din_a[46] & din_b[42]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_49  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[42]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_47_sumout ),
	.cout(Xd_0__inst_mult_3_48 ),
	.shareout(Xd_0__inst_mult_3_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_116 (
// Equation(s):
// Xd_0__inst_mult_0_364  = SUM(( !Xd_0__inst_mult_0_552  $ (!Xd_0__inst_mult_0_556 ) ) + ( Xd_0__inst_mult_0_358  ) + ( Xd_0__inst_mult_0_357  ))
// Xd_0__inst_mult_0_365  = CARRY(( !Xd_0__inst_mult_0_552  $ (!Xd_0__inst_mult_0_556 ) ) + ( Xd_0__inst_mult_0_358  ) + ( Xd_0__inst_mult_0_357  ))
// Xd_0__inst_mult_0_366  = SHARE((Xd_0__inst_mult_0_552  & Xd_0__inst_mult_0_556 ))

	.dataa(!Xd_0__inst_mult_0_552 ),
	.datab(!Xd_0__inst_mult_0_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_357 ),
	.sharein(Xd_0__inst_mult_0_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_364 ),
	.cout(Xd_0__inst_mult_0_365 ),
	.shareout(Xd_0__inst_mult_0_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_39 (
// Equation(s):
// Xd_0__inst_mult_0_39_sumout  = SUM(( (din_a[10] & din_b[6]) ) + ( Xd_0__inst_mult_1_45  ) + ( Xd_0__inst_mult_1_44  ))
// Xd_0__inst_mult_0_40  = CARRY(( (din_a[10] & din_b[6]) ) + ( Xd_0__inst_mult_1_45  ) + ( Xd_0__inst_mult_1_44  ))
// Xd_0__inst_mult_0_41  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_44 ),
	.sharein(Xd_0__inst_mult_1_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_39_sumout ),
	.cout(Xd_0__inst_mult_0_40 ),
	.shareout(Xd_0__inst_mult_0_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_116 (
// Equation(s):
// Xd_0__inst_mult_1_364  = SUM(( !Xd_0__inst_mult_1_556  $ (!Xd_0__inst_mult_1_560 ) ) + ( Xd_0__inst_mult_1_358  ) + ( Xd_0__inst_mult_1_357  ))
// Xd_0__inst_mult_1_365  = CARRY(( !Xd_0__inst_mult_1_556  $ (!Xd_0__inst_mult_1_560 ) ) + ( Xd_0__inst_mult_1_358  ) + ( Xd_0__inst_mult_1_357  ))
// Xd_0__inst_mult_1_366  = SHARE((Xd_0__inst_mult_1_556  & Xd_0__inst_mult_1_560 ))

	.dataa(!Xd_0__inst_mult_1_556 ),
	.datab(!Xd_0__inst_mult_1_560 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_357 ),
	.sharein(Xd_0__inst_mult_1_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_364 ),
	.cout(Xd_0__inst_mult_1_365 ),
	.shareout(Xd_0__inst_mult_1_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_43 (
// Equation(s):
// Xd_0__inst_mult_1_43_sumout  = SUM(( (din_a[22] & din_b[18]) ) + ( Xd_0__inst_mult_14_57  ) + ( Xd_0__inst_mult_14_56  ))
// Xd_0__inst_mult_1_44  = CARRY(( (din_a[22] & din_b[18]) ) + ( Xd_0__inst_mult_14_57  ) + ( Xd_0__inst_mult_14_56  ))
// Xd_0__inst_mult_1_45  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_56 ),
	.sharein(Xd_0__inst_mult_14_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_43_sumout ),
	.cout(Xd_0__inst_mult_1_44 ),
	.shareout(Xd_0__inst_mult_1_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_120 (
// Equation(s):
// Xd_0__inst_mult_12_392  = SUM(( !Xd_0__inst_mult_12_564  $ (!Xd_0__inst_mult_12_180  $ (((din_a[153] & din_b[152])))) ) + ( Xd_0__inst_mult_12_390  ) + ( Xd_0__inst_mult_12_389  ))
// Xd_0__inst_mult_12_393  = CARRY(( !Xd_0__inst_mult_12_564  $ (!Xd_0__inst_mult_12_180  $ (((din_a[153] & din_b[152])))) ) + ( Xd_0__inst_mult_12_390  ) + ( Xd_0__inst_mult_12_389  ))
// Xd_0__inst_mult_12_394  = SHARE((!Xd_0__inst_mult_12_564  & (Xd_0__inst_mult_12_180  & (din_a[153] & din_b[152]))) # (Xd_0__inst_mult_12_564  & (((din_a[153] & din_b[152])) # (Xd_0__inst_mult_12_180 ))))

	.dataa(!Xd_0__inst_mult_12_564 ),
	.datab(!Xd_0__inst_mult_12_180 ),
	.datac(!din_a[153]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_389 ),
	.sharein(Xd_0__inst_mult_12_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_392 ),
	.cout(Xd_0__inst_mult_12_393 ),
	.shareout(Xd_0__inst_mult_12_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_51 (
// Equation(s):
// Xd_0__inst_mult_12_51_sumout  = SUM(( (din_a[154] & din_b[151]) ) + ( Xd_0__inst_mult_13_49  ) + ( Xd_0__inst_mult_13_48  ))
// Xd_0__inst_mult_12_52  = CARRY(( (din_a[154] & din_b[151]) ) + ( Xd_0__inst_mult_13_49  ) + ( Xd_0__inst_mult_13_48  ))
// Xd_0__inst_mult_12_53  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_48 ),
	.sharein(Xd_0__inst_mult_13_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_51_sumout ),
	.cout(Xd_0__inst_mult_12_52 ),
	.shareout(Xd_0__inst_mult_12_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_118 (
// Equation(s):
// Xd_0__inst_mult_13_372  = SUM(( !Xd_0__inst_mult_13_560  $ (!Xd_0__inst_mult_13_564  $ (((din_a[165] & din_b[164])))) ) + ( Xd_0__inst_mult_13_370  ) + ( Xd_0__inst_mult_13_369  ))
// Xd_0__inst_mult_13_373  = CARRY(( !Xd_0__inst_mult_13_560  $ (!Xd_0__inst_mult_13_564  $ (((din_a[165] & din_b[164])))) ) + ( Xd_0__inst_mult_13_370  ) + ( Xd_0__inst_mult_13_369  ))
// Xd_0__inst_mult_13_374  = SHARE((!Xd_0__inst_mult_13_560  & (Xd_0__inst_mult_13_564  & (din_a[165] & din_b[164]))) # (Xd_0__inst_mult_13_560  & (((din_a[165] & din_b[164])) # (Xd_0__inst_mult_13_564 ))))

	.dataa(!Xd_0__inst_mult_13_560 ),
	.datab(!Xd_0__inst_mult_13_564 ),
	.datac(!din_a[165]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_369 ),
	.sharein(Xd_0__inst_mult_13_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_372 ),
	.cout(Xd_0__inst_mult_13_373 ),
	.shareout(Xd_0__inst_mult_13_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_47 (
// Equation(s):
// Xd_0__inst_mult_13_47_sumout  = SUM(( (din_a[166] & din_b[163]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_48  = CARRY(( (din_a[166] & din_b[163]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_49  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[163]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_13_47_sumout ),
	.cout(Xd_0__inst_mult_13_48 ),
	.shareout(Xd_0__inst_mult_13_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_122 (
// Equation(s):
// Xd_0__inst_mult_14_388  = SUM(( !Xd_0__inst_mult_14_564  $ (!Xd_0__inst_mult_14_568  $ (((din_a[177] & din_b[176])))) ) + ( Xd_0__inst_mult_14_386  ) + ( Xd_0__inst_mult_14_385  ))
// Xd_0__inst_mult_14_389  = CARRY(( !Xd_0__inst_mult_14_564  $ (!Xd_0__inst_mult_14_568  $ (((din_a[177] & din_b[176])))) ) + ( Xd_0__inst_mult_14_386  ) + ( Xd_0__inst_mult_14_385  ))
// Xd_0__inst_mult_14_390  = SHARE((!Xd_0__inst_mult_14_564  & (Xd_0__inst_mult_14_568  & (din_a[177] & din_b[176]))) # (Xd_0__inst_mult_14_564  & (((din_a[177] & din_b[176])) # (Xd_0__inst_mult_14_568 ))))

	.dataa(!Xd_0__inst_mult_14_564 ),
	.datab(!Xd_0__inst_mult_14_568 ),
	.datac(!din_a[177]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_385 ),
	.sharein(Xd_0__inst_mult_14_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_388 ),
	.cout(Xd_0__inst_mult_14_389 ),
	.shareout(Xd_0__inst_mult_14_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_55 (
// Equation(s):
// Xd_0__inst_mult_14_55_sumout  = SUM(( (din_a[178] & din_b[175]) ) + ( Xd_0__inst_mult_15_53  ) + ( Xd_0__inst_mult_15_52  ))
// Xd_0__inst_mult_14_56  = CARRY(( (din_a[178] & din_b[175]) ) + ( Xd_0__inst_mult_15_53  ) + ( Xd_0__inst_mult_15_52  ))
// Xd_0__inst_mult_14_57  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[175]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_52 ),
	.sharein(Xd_0__inst_mult_15_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_55_sumout ),
	.cout(Xd_0__inst_mult_14_56 ),
	.shareout(Xd_0__inst_mult_14_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_124 (
// Equation(s):
// Xd_0__inst_mult_15_396  = SUM(( !Xd_0__inst_mult_15_572  $ (!Xd_0__inst_mult_15_180  $ (((din_a[189] & din_b[188])))) ) + ( Xd_0__inst_mult_15_394  ) + ( Xd_0__inst_mult_15_393  ))
// Xd_0__inst_mult_15_397  = CARRY(( !Xd_0__inst_mult_15_572  $ (!Xd_0__inst_mult_15_180  $ (((din_a[189] & din_b[188])))) ) + ( Xd_0__inst_mult_15_394  ) + ( Xd_0__inst_mult_15_393  ))
// Xd_0__inst_mult_15_398  = SHARE((!Xd_0__inst_mult_15_572  & (Xd_0__inst_mult_15_180  & (din_a[189] & din_b[188]))) # (Xd_0__inst_mult_15_572  & (((din_a[189] & din_b[188])) # (Xd_0__inst_mult_15_180 ))))

	.dataa(!Xd_0__inst_mult_15_572 ),
	.datab(!Xd_0__inst_mult_15_180 ),
	.datac(!din_a[189]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_393 ),
	.sharein(Xd_0__inst_mult_15_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_396 ),
	.cout(Xd_0__inst_mult_15_397 ),
	.shareout(Xd_0__inst_mult_15_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_51 (
// Equation(s):
// Xd_0__inst_mult_15_51_sumout  = SUM(( (din_a[190] & din_b[187]) ) + ( Xd_0__inst_mult_12_53  ) + ( Xd_0__inst_mult_12_52  ))
// Xd_0__inst_mult_15_52  = CARRY(( (din_a[190] & din_b[187]) ) + ( Xd_0__inst_mult_12_53  ) + ( Xd_0__inst_mult_12_52  ))
// Xd_0__inst_mult_15_53  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[187]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_52 ),
	.sharein(Xd_0__inst_mult_12_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_51_sumout ),
	.cout(Xd_0__inst_mult_15_52 ),
	.shareout(Xd_0__inst_mult_15_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_114 (
// Equation(s):
// Xd_0__inst_mult_10_368  = SUM(( !Xd_0__inst_mult_10_556  $ (!Xd_0__inst_mult_10_560  $ (((din_a[129] & din_b[128])))) ) + ( Xd_0__inst_mult_10_366  ) + ( Xd_0__inst_mult_10_365  ))
// Xd_0__inst_mult_10_369  = CARRY(( !Xd_0__inst_mult_10_556  $ (!Xd_0__inst_mult_10_560  $ (((din_a[129] & din_b[128])))) ) + ( Xd_0__inst_mult_10_366  ) + ( Xd_0__inst_mult_10_365  ))
// Xd_0__inst_mult_10_370  = SHARE((!Xd_0__inst_mult_10_556  & (Xd_0__inst_mult_10_560  & (din_a[129] & din_b[128]))) # (Xd_0__inst_mult_10_556  & (((din_a[129] & din_b[128])) # (Xd_0__inst_mult_10_560 ))))

	.dataa(!Xd_0__inst_mult_10_556 ),
	.datab(!Xd_0__inst_mult_10_560 ),
	.datac(!din_a[129]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_365 ),
	.sharein(Xd_0__inst_mult_10_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_368 ),
	.cout(Xd_0__inst_mult_10_369 ),
	.shareout(Xd_0__inst_mult_10_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_43 (
// Equation(s):
// Xd_0__inst_mult_10_43_sumout  = SUM(( (din_a[130] & din_b[127]) ) + ( Xd_0__inst_mult_11_45  ) + ( Xd_0__inst_mult_11_44  ))
// Xd_0__inst_mult_10_44  = CARRY(( (din_a[130] & din_b[127]) ) + ( Xd_0__inst_mult_11_45  ) + ( Xd_0__inst_mult_11_44  ))
// Xd_0__inst_mult_10_45  = SHARE(GND)

	.dataa(!din_a[130]),
	.datab(!din_b[127]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_44 ),
	.sharein(Xd_0__inst_mult_11_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_43_sumout ),
	.cout(Xd_0__inst_mult_10_44 ),
	.shareout(Xd_0__inst_mult_10_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_118 (
// Equation(s):
// Xd_0__inst_mult_11_372  = SUM(( !Xd_0__inst_mult_11_560  $ (!Xd_0__inst_mult_11_564  $ (((din_a[141] & din_b[140])))) ) + ( Xd_0__inst_mult_11_370  ) + ( Xd_0__inst_mult_11_369  ))
// Xd_0__inst_mult_11_373  = CARRY(( !Xd_0__inst_mult_11_560  $ (!Xd_0__inst_mult_11_564  $ (((din_a[141] & din_b[140])))) ) + ( Xd_0__inst_mult_11_370  ) + ( Xd_0__inst_mult_11_369  ))
// Xd_0__inst_mult_11_374  = SHARE((!Xd_0__inst_mult_11_560  & (Xd_0__inst_mult_11_564  & (din_a[141] & din_b[140]))) # (Xd_0__inst_mult_11_560  & (((din_a[141] & din_b[140])) # (Xd_0__inst_mult_11_564 ))))

	.dataa(!Xd_0__inst_mult_11_560 ),
	.datab(!Xd_0__inst_mult_11_564 ),
	.datac(!din_a[141]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_369 ),
	.sharein(Xd_0__inst_mult_11_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_372 ),
	.cout(Xd_0__inst_mult_11_373 ),
	.shareout(Xd_0__inst_mult_11_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_43 (
// Equation(s):
// Xd_0__inst_mult_11_43_sumout  = SUM(( (din_a[142] & din_b[139]) ) + ( Xd_0__inst_mult_8_53  ) + ( Xd_0__inst_mult_8_52  ))
// Xd_0__inst_mult_11_44  = CARRY(( (din_a[142] & din_b[139]) ) + ( Xd_0__inst_mult_8_53  ) + ( Xd_0__inst_mult_8_52  ))
// Xd_0__inst_mult_11_45  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[139]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_52 ),
	.sharein(Xd_0__inst_mult_8_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_43_sumout ),
	.cout(Xd_0__inst_mult_11_44 ),
	.shareout(Xd_0__inst_mult_11_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_118 (
// Equation(s):
// Xd_0__inst_mult_8_372  = SUM(( !Xd_0__inst_mult_8_560  $ (!Xd_0__inst_mult_8_564  $ (((din_a[105] & din_b[104])))) ) + ( Xd_0__inst_mult_8_370  ) + ( Xd_0__inst_mult_8_369  ))
// Xd_0__inst_mult_8_373  = CARRY(( !Xd_0__inst_mult_8_560  $ (!Xd_0__inst_mult_8_564  $ (((din_a[105] & din_b[104])))) ) + ( Xd_0__inst_mult_8_370  ) + ( Xd_0__inst_mult_8_369  ))
// Xd_0__inst_mult_8_374  = SHARE((!Xd_0__inst_mult_8_560  & (Xd_0__inst_mult_8_564  & (din_a[105] & din_b[104]))) # (Xd_0__inst_mult_8_560  & (((din_a[105] & din_b[104])) # (Xd_0__inst_mult_8_564 ))))

	.dataa(!Xd_0__inst_mult_8_560 ),
	.datab(!Xd_0__inst_mult_8_564 ),
	.datac(!din_a[105]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_369 ),
	.sharein(Xd_0__inst_mult_8_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_372 ),
	.cout(Xd_0__inst_mult_8_373 ),
	.shareout(Xd_0__inst_mult_8_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_51 (
// Equation(s):
// Xd_0__inst_mult_8_51_sumout  = SUM(( (din_a[106] & din_b[103]) ) + ( Xd_0__inst_i29_27  ) + ( Xd_0__inst_i29_26  ))
// Xd_0__inst_mult_8_52  = CARRY(( (din_a[106] & din_b[103]) ) + ( Xd_0__inst_i29_27  ) + ( Xd_0__inst_i29_26  ))
// Xd_0__inst_mult_8_53  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_26 ),
	.sharein(Xd_0__inst_i29_27 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_51_sumout ),
	.cout(Xd_0__inst_mult_8_52 ),
	.shareout(Xd_0__inst_mult_8_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_114 (
// Equation(s):
// Xd_0__inst_mult_9_368  = SUM(( !Xd_0__inst_mult_9_556  $ (!Xd_0__inst_mult_9_560  $ (((din_a[117] & din_b[116])))) ) + ( Xd_0__inst_mult_9_366  ) + ( Xd_0__inst_mult_9_365  ))
// Xd_0__inst_mult_9_369  = CARRY(( !Xd_0__inst_mult_9_556  $ (!Xd_0__inst_mult_9_560  $ (((din_a[117] & din_b[116])))) ) + ( Xd_0__inst_mult_9_366  ) + ( Xd_0__inst_mult_9_365  ))
// Xd_0__inst_mult_9_370  = SHARE((!Xd_0__inst_mult_9_556  & (Xd_0__inst_mult_9_560  & (din_a[117] & din_b[116]))) # (Xd_0__inst_mult_9_556  & (((din_a[117] & din_b[116])) # (Xd_0__inst_mult_9_560 ))))

	.dataa(!Xd_0__inst_mult_9_556 ),
	.datab(!Xd_0__inst_mult_9_560 ),
	.datac(!din_a[117]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_365 ),
	.sharein(Xd_0__inst_mult_9_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_368 ),
	.cout(Xd_0__inst_mult_9_369 ),
	.shareout(Xd_0__inst_mult_9_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_114 (
// Equation(s):
// Xd_0__inst_mult_6_368  = SUM(( !Xd_0__inst_mult_6_556  $ (!Xd_0__inst_mult_6_560  $ (((din_a[81] & din_b[80])))) ) + ( Xd_0__inst_mult_6_366  ) + ( Xd_0__inst_mult_6_365  ))
// Xd_0__inst_mult_6_369  = CARRY(( !Xd_0__inst_mult_6_556  $ (!Xd_0__inst_mult_6_560  $ (((din_a[81] & din_b[80])))) ) + ( Xd_0__inst_mult_6_366  ) + ( Xd_0__inst_mult_6_365  ))
// Xd_0__inst_mult_6_370  = SHARE((!Xd_0__inst_mult_6_556  & (Xd_0__inst_mult_6_560  & (din_a[81] & din_b[80]))) # (Xd_0__inst_mult_6_556  & (((din_a[81] & din_b[80])) # (Xd_0__inst_mult_6_560 ))))

	.dataa(!Xd_0__inst_mult_6_556 ),
	.datab(!Xd_0__inst_mult_6_560 ),
	.datac(!din_a[81]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_365 ),
	.sharein(Xd_0__inst_mult_6_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_368 ),
	.cout(Xd_0__inst_mult_6_369 ),
	.shareout(Xd_0__inst_mult_6_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_47 (
// Equation(s):
// Xd_0__inst_mult_6_47_sumout  = SUM(( (din_a[82] & din_b[79]) ) + ( Xd_0__inst_mult_7_41  ) + ( Xd_0__inst_mult_7_40  ))
// Xd_0__inst_mult_6_48  = CARRY(( (din_a[82] & din_b[79]) ) + ( Xd_0__inst_mult_7_41  ) + ( Xd_0__inst_mult_7_40  ))
// Xd_0__inst_mult_6_49  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_40 ),
	.sharein(Xd_0__inst_mult_7_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_47_sumout ),
	.cout(Xd_0__inst_mult_6_48 ),
	.shareout(Xd_0__inst_mult_6_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_112 (
// Equation(s):
// Xd_0__inst_mult_7_360  = SUM(( !Xd_0__inst_mult_7_556  $ (!Xd_0__inst_mult_7_560  $ (((din_a[93] & din_b[92])))) ) + ( Xd_0__inst_mult_7_358  ) + ( Xd_0__inst_mult_7_357  ))
// Xd_0__inst_mult_7_361  = CARRY(( !Xd_0__inst_mult_7_556  $ (!Xd_0__inst_mult_7_560  $ (((din_a[93] & din_b[92])))) ) + ( Xd_0__inst_mult_7_358  ) + ( Xd_0__inst_mult_7_357  ))
// Xd_0__inst_mult_7_362  = SHARE((!Xd_0__inst_mult_7_556  & (Xd_0__inst_mult_7_560  & (din_a[93] & din_b[92]))) # (Xd_0__inst_mult_7_556  & (((din_a[93] & din_b[92])) # (Xd_0__inst_mult_7_560 ))))

	.dataa(!Xd_0__inst_mult_7_556 ),
	.datab(!Xd_0__inst_mult_7_560 ),
	.datac(!din_a[93]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_357 ),
	.sharein(Xd_0__inst_mult_7_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_360 ),
	.cout(Xd_0__inst_mult_7_361 ),
	.shareout(Xd_0__inst_mult_7_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_39 (
// Equation(s):
// Xd_0__inst_mult_7_39_sumout  = SUM(( (din_a[94] & din_b[91]) ) + ( Xd_0__inst_mult_4_45  ) + ( Xd_0__inst_mult_4_44  ))
// Xd_0__inst_mult_7_40  = CARRY(( (din_a[94] & din_b[91]) ) + ( Xd_0__inst_mult_4_45  ) + ( Xd_0__inst_mult_4_44  ))
// Xd_0__inst_mult_7_41  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_44 ),
	.sharein(Xd_0__inst_mult_4_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_39_sumout ),
	.cout(Xd_0__inst_mult_7_40 ),
	.shareout(Xd_0__inst_mult_7_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_124 (
// Equation(s):
// Xd_0__inst_mult_4_396  = SUM(( !Xd_0__inst_mult_4_568  $ (!Xd_0__inst_mult_4_180  $ (((din_a[57] & din_b[56])))) ) + ( Xd_0__inst_mult_4_394  ) + ( Xd_0__inst_mult_4_393  ))
// Xd_0__inst_mult_4_397  = CARRY(( !Xd_0__inst_mult_4_568  $ (!Xd_0__inst_mult_4_180  $ (((din_a[57] & din_b[56])))) ) + ( Xd_0__inst_mult_4_394  ) + ( Xd_0__inst_mult_4_393  ))
// Xd_0__inst_mult_4_398  = SHARE((!Xd_0__inst_mult_4_568  & (Xd_0__inst_mult_4_180  & (din_a[57] & din_b[56]))) # (Xd_0__inst_mult_4_568  & (((din_a[57] & din_b[56])) # (Xd_0__inst_mult_4_180 ))))

	.dataa(!Xd_0__inst_mult_4_568 ),
	.datab(!Xd_0__inst_mult_4_180 ),
	.datac(!din_a[57]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_393 ),
	.sharein(Xd_0__inst_mult_4_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_396 ),
	.cout(Xd_0__inst_mult_4_397 ),
	.shareout(Xd_0__inst_mult_4_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_43 (
// Equation(s):
// Xd_0__inst_mult_4_43_sumout  = SUM(( (din_a[58] & din_b[55]) ) + ( Xd_0__inst_mult_5_49  ) + ( Xd_0__inst_mult_5_48  ))
// Xd_0__inst_mult_4_44  = CARRY(( (din_a[58] & din_b[55]) ) + ( Xd_0__inst_mult_5_49  ) + ( Xd_0__inst_mult_5_48  ))
// Xd_0__inst_mult_4_45  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_48 ),
	.sharein(Xd_0__inst_mult_5_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_43_sumout ),
	.cout(Xd_0__inst_mult_4_44 ),
	.shareout(Xd_0__inst_mult_4_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_112 (
// Equation(s):
// Xd_0__inst_mult_5_360  = SUM(( !Xd_0__inst_mult_5_556  $ (!Xd_0__inst_mult_5_560  $ (((din_a[69] & din_b[68])))) ) + ( Xd_0__inst_mult_5_358  ) + ( Xd_0__inst_mult_5_357  ))
// Xd_0__inst_mult_5_361  = CARRY(( !Xd_0__inst_mult_5_556  $ (!Xd_0__inst_mult_5_560  $ (((din_a[69] & din_b[68])))) ) + ( Xd_0__inst_mult_5_358  ) + ( Xd_0__inst_mult_5_357  ))
// Xd_0__inst_mult_5_362  = SHARE((!Xd_0__inst_mult_5_556  & (Xd_0__inst_mult_5_560  & (din_a[69] & din_b[68]))) # (Xd_0__inst_mult_5_556  & (((din_a[69] & din_b[68])) # (Xd_0__inst_mult_5_560 ))))

	.dataa(!Xd_0__inst_mult_5_556 ),
	.datab(!Xd_0__inst_mult_5_560 ),
	.datac(!din_a[69]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_357 ),
	.sharein(Xd_0__inst_mult_5_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_360 ),
	.cout(Xd_0__inst_mult_5_361 ),
	.shareout(Xd_0__inst_mult_5_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_47 (
// Equation(s):
// Xd_0__inst_mult_5_47_sumout  = SUM(( (din_a[70] & din_b[67]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_48  = CARRY(( (din_a[70] & din_b[67]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_49  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_47_sumout ),
	.cout(Xd_0__inst_mult_5_48 ),
	.shareout(Xd_0__inst_mult_5_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_116 (
// Equation(s):
// Xd_0__inst_mult_2_364  = SUM(( !Xd_0__inst_mult_2_560  $ (!Xd_0__inst_mult_2_564  $ (((din_a[33] & din_b[32])))) ) + ( Xd_0__inst_mult_2_362  ) + ( Xd_0__inst_mult_2_361  ))
// Xd_0__inst_mult_2_365  = CARRY(( !Xd_0__inst_mult_2_560  $ (!Xd_0__inst_mult_2_564  $ (((din_a[33] & din_b[32])))) ) + ( Xd_0__inst_mult_2_362  ) + ( Xd_0__inst_mult_2_361  ))
// Xd_0__inst_mult_2_366  = SHARE((!Xd_0__inst_mult_2_560  & (Xd_0__inst_mult_2_564  & (din_a[33] & din_b[32]))) # (Xd_0__inst_mult_2_560  & (((din_a[33] & din_b[32])) # (Xd_0__inst_mult_2_564 ))))

	.dataa(!Xd_0__inst_mult_2_560 ),
	.datab(!Xd_0__inst_mult_2_564 ),
	.datac(!din_a[33]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_361 ),
	.sharein(Xd_0__inst_mult_2_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_364 ),
	.cout(Xd_0__inst_mult_2_365 ),
	.shareout(Xd_0__inst_mult_2_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_47 (
// Equation(s):
// Xd_0__inst_mult_2_47_sumout  = SUM(( (din_a[34] & din_b[31]) ) + ( Xd_0__inst_mult_3_53  ) + ( Xd_0__inst_mult_3_52  ))
// Xd_0__inst_mult_2_48  = CARRY(( (din_a[34] & din_b[31]) ) + ( Xd_0__inst_mult_3_53  ) + ( Xd_0__inst_mult_3_52  ))
// Xd_0__inst_mult_2_49  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_52 ),
	.sharein(Xd_0__inst_mult_3_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_47_sumout ),
	.cout(Xd_0__inst_mult_2_48 ),
	.shareout(Xd_0__inst_mult_2_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_112 (
// Equation(s):
// Xd_0__inst_mult_3_360  = SUM(( !Xd_0__inst_mult_3_556  $ (!Xd_0__inst_mult_3_560  $ (((din_a[45] & din_b[44])))) ) + ( Xd_0__inst_mult_3_358  ) + ( Xd_0__inst_mult_3_357  ))
// Xd_0__inst_mult_3_361  = CARRY(( !Xd_0__inst_mult_3_556  $ (!Xd_0__inst_mult_3_560  $ (((din_a[45] & din_b[44])))) ) + ( Xd_0__inst_mult_3_358  ) + ( Xd_0__inst_mult_3_357  ))
// Xd_0__inst_mult_3_362  = SHARE((!Xd_0__inst_mult_3_556  & (Xd_0__inst_mult_3_560  & (din_a[45] & din_b[44]))) # (Xd_0__inst_mult_3_556  & (((din_a[45] & din_b[44])) # (Xd_0__inst_mult_3_560 ))))

	.dataa(!Xd_0__inst_mult_3_556 ),
	.datab(!Xd_0__inst_mult_3_560 ),
	.datac(!din_a[45]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_357 ),
	.sharein(Xd_0__inst_mult_3_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_360 ),
	.cout(Xd_0__inst_mult_3_361 ),
	.shareout(Xd_0__inst_mult_3_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_51 (
// Equation(s):
// Xd_0__inst_mult_3_51_sumout  = SUM(( (din_a[46] & din_b[43]) ) + ( Xd_0__inst_mult_0_45  ) + ( Xd_0__inst_mult_0_44  ))
// Xd_0__inst_mult_3_52  = CARRY(( (din_a[46] & din_b[43]) ) + ( Xd_0__inst_mult_0_45  ) + ( Xd_0__inst_mult_0_44  ))
// Xd_0__inst_mult_3_53  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_44 ),
	.sharein(Xd_0__inst_mult_0_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_51_sumout ),
	.cout(Xd_0__inst_mult_3_52 ),
	.shareout(Xd_0__inst_mult_3_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_117 (
// Equation(s):
// Xd_0__inst_mult_0_368  = SUM(( !Xd_0__inst_mult_0_560  $ (!Xd_0__inst_mult_0_564  $ (((din_a[9] & din_b[8])))) ) + ( Xd_0__inst_mult_0_366  ) + ( Xd_0__inst_mult_0_365  ))
// Xd_0__inst_mult_0_369  = CARRY(( !Xd_0__inst_mult_0_560  $ (!Xd_0__inst_mult_0_564  $ (((din_a[9] & din_b[8])))) ) + ( Xd_0__inst_mult_0_366  ) + ( Xd_0__inst_mult_0_365  ))
// Xd_0__inst_mult_0_370  = SHARE((!Xd_0__inst_mult_0_560  & (Xd_0__inst_mult_0_564  & (din_a[9] & din_b[8]))) # (Xd_0__inst_mult_0_560  & (((din_a[9] & din_b[8])) # (Xd_0__inst_mult_0_564 ))))

	.dataa(!Xd_0__inst_mult_0_560 ),
	.datab(!Xd_0__inst_mult_0_564 ),
	.datac(!din_a[9]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_365 ),
	.sharein(Xd_0__inst_mult_0_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_368 ),
	.cout(Xd_0__inst_mult_0_369 ),
	.shareout(Xd_0__inst_mult_0_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_43 (
// Equation(s):
// Xd_0__inst_mult_0_43_sumout  = SUM(( (din_a[10] & din_b[7]) ) + ( Xd_0__inst_mult_1_49  ) + ( Xd_0__inst_mult_1_48  ))
// Xd_0__inst_mult_0_44  = CARRY(( (din_a[10] & din_b[7]) ) + ( Xd_0__inst_mult_1_49  ) + ( Xd_0__inst_mult_1_48  ))
// Xd_0__inst_mult_0_45  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_48 ),
	.sharein(Xd_0__inst_mult_1_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_43_sumout ),
	.cout(Xd_0__inst_mult_0_44 ),
	.shareout(Xd_0__inst_mult_0_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_117 (
// Equation(s):
// Xd_0__inst_mult_1_368  = SUM(( !Xd_0__inst_mult_1_564  $ (!Xd_0__inst_mult_1_568  $ (((din_a[21] & din_b[20])))) ) + ( Xd_0__inst_mult_1_366  ) + ( Xd_0__inst_mult_1_365  ))
// Xd_0__inst_mult_1_369  = CARRY(( !Xd_0__inst_mult_1_564  $ (!Xd_0__inst_mult_1_568  $ (((din_a[21] & din_b[20])))) ) + ( Xd_0__inst_mult_1_366  ) + ( Xd_0__inst_mult_1_365  ))
// Xd_0__inst_mult_1_370  = SHARE((!Xd_0__inst_mult_1_564  & (Xd_0__inst_mult_1_568  & (din_a[21] & din_b[20]))) # (Xd_0__inst_mult_1_564  & (((din_a[21] & din_b[20])) # (Xd_0__inst_mult_1_568 ))))

	.dataa(!Xd_0__inst_mult_1_564 ),
	.datab(!Xd_0__inst_mult_1_568 ),
	.datac(!din_a[21]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_365 ),
	.sharein(Xd_0__inst_mult_1_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_368 ),
	.cout(Xd_0__inst_mult_1_369 ),
	.shareout(Xd_0__inst_mult_1_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_47 (
// Equation(s):
// Xd_0__inst_mult_1_47_sumout  = SUM(( (din_a[22] & din_b[19]) ) + ( Xd_0__inst_mult_14_61  ) + ( Xd_0__inst_mult_14_60  ))
// Xd_0__inst_mult_1_48  = CARRY(( (din_a[22] & din_b[19]) ) + ( Xd_0__inst_mult_14_61  ) + ( Xd_0__inst_mult_14_60  ))
// Xd_0__inst_mult_1_49  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_60 ),
	.sharein(Xd_0__inst_mult_14_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_47_sumout ),
	.cout(Xd_0__inst_mult_1_48 ),
	.shareout(Xd_0__inst_mult_1_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_121 (
// Equation(s):
// Xd_0__inst_mult_12_396  = SUM(( !Xd_0__inst_mult_12_173  $ (((!din_a[153]) # (!din_b[153]))) ) + ( Xd_0__inst_mult_12_394  ) + ( Xd_0__inst_mult_12_393  ))
// Xd_0__inst_mult_12_397  = CARRY(( !Xd_0__inst_mult_12_173  $ (((!din_a[153]) # (!din_b[153]))) ) + ( Xd_0__inst_mult_12_394  ) + ( Xd_0__inst_mult_12_393  ))
// Xd_0__inst_mult_12_398  = SHARE((din_a[153] & (din_b[153] & Xd_0__inst_mult_12_173 )))

	.dataa(!din_a[153]),
	.datab(!din_b[153]),
	.datac(!Xd_0__inst_mult_12_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_393 ),
	.sharein(Xd_0__inst_mult_12_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_396 ),
	.cout(Xd_0__inst_mult_12_397 ),
	.shareout(Xd_0__inst_mult_12_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_55 (
// Equation(s):
// Xd_0__inst_mult_12_55_sumout  = SUM(( (din_a[154] & din_b[152]) ) + ( Xd_0__inst_mult_13_53  ) + ( Xd_0__inst_mult_13_52  ))
// Xd_0__inst_mult_12_56  = CARRY(( (din_a[154] & din_b[152]) ) + ( Xd_0__inst_mult_13_53  ) + ( Xd_0__inst_mult_13_52  ))
// Xd_0__inst_mult_12_57  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[152]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_52 ),
	.sharein(Xd_0__inst_mult_13_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_55_sumout ),
	.cout(Xd_0__inst_mult_12_56 ),
	.shareout(Xd_0__inst_mult_12_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_119 (
// Equation(s):
// Xd_0__inst_mult_13_376  = SUM(( !Xd_0__inst_mult_13_568  $ (((!din_a[165]) # (!din_b[165]))) ) + ( Xd_0__inst_mult_13_374  ) + ( Xd_0__inst_mult_13_373  ))
// Xd_0__inst_mult_13_377  = CARRY(( !Xd_0__inst_mult_13_568  $ (((!din_a[165]) # (!din_b[165]))) ) + ( Xd_0__inst_mult_13_374  ) + ( Xd_0__inst_mult_13_373  ))
// Xd_0__inst_mult_13_378  = SHARE((din_a[165] & (din_b[165] & Xd_0__inst_mult_13_568 )))

	.dataa(!din_a[165]),
	.datab(!din_b[165]),
	.datac(!Xd_0__inst_mult_13_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_373 ),
	.sharein(Xd_0__inst_mult_13_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_376 ),
	.cout(Xd_0__inst_mult_13_377 ),
	.shareout(Xd_0__inst_mult_13_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_51 (
// Equation(s):
// Xd_0__inst_mult_13_51_sumout  = SUM(( (din_a[166] & din_b[164]) ) + ( Xd_0__inst_mult_10_49  ) + ( Xd_0__inst_mult_10_48  ))
// Xd_0__inst_mult_13_52  = CARRY(( (din_a[166] & din_b[164]) ) + ( Xd_0__inst_mult_10_49  ) + ( Xd_0__inst_mult_10_48  ))
// Xd_0__inst_mult_13_53  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[164]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_48 ),
	.sharein(Xd_0__inst_mult_10_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_51_sumout ),
	.cout(Xd_0__inst_mult_13_52 ),
	.shareout(Xd_0__inst_mult_13_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_123 (
// Equation(s):
// Xd_0__inst_mult_14_392  = SUM(( !Xd_0__inst_mult_14_572  $ (((!din_a[177]) # (!din_b[177]))) ) + ( Xd_0__inst_mult_14_390  ) + ( Xd_0__inst_mult_14_389  ))
// Xd_0__inst_mult_14_393  = CARRY(( !Xd_0__inst_mult_14_572  $ (((!din_a[177]) # (!din_b[177]))) ) + ( Xd_0__inst_mult_14_390  ) + ( Xd_0__inst_mult_14_389  ))
// Xd_0__inst_mult_14_394  = SHARE((din_a[177] & (din_b[177] & Xd_0__inst_mult_14_572 )))

	.dataa(!din_a[177]),
	.datab(!din_b[177]),
	.datac(!Xd_0__inst_mult_14_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_389 ),
	.sharein(Xd_0__inst_mult_14_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_392 ),
	.cout(Xd_0__inst_mult_14_393 ),
	.shareout(Xd_0__inst_mult_14_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_59 (
// Equation(s):
// Xd_0__inst_mult_14_59_sumout  = SUM(( (din_a[178] & din_b[176]) ) + ( Xd_0__inst_mult_1_57  ) + ( Xd_0__inst_mult_1_56  ))
// Xd_0__inst_mult_14_60  = CARRY(( (din_a[178] & din_b[176]) ) + ( Xd_0__inst_mult_1_57  ) + ( Xd_0__inst_mult_1_56  ))
// Xd_0__inst_mult_14_61  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[176]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_56 ),
	.sharein(Xd_0__inst_mult_1_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_59_sumout ),
	.cout(Xd_0__inst_mult_14_60 ),
	.shareout(Xd_0__inst_mult_14_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_125 (
// Equation(s):
// Xd_0__inst_mult_15_400  = SUM(( !Xd_0__inst_mult_15_177  $ (((!din_a[189]) # (!din_b[189]))) ) + ( Xd_0__inst_mult_15_398  ) + ( Xd_0__inst_mult_15_397  ))
// Xd_0__inst_mult_15_401  = CARRY(( !Xd_0__inst_mult_15_177  $ (((!din_a[189]) # (!din_b[189]))) ) + ( Xd_0__inst_mult_15_398  ) + ( Xd_0__inst_mult_15_397  ))
// Xd_0__inst_mult_15_402  = SHARE((din_a[189] & (din_b[189] & Xd_0__inst_mult_15_177 )))

	.dataa(!din_a[189]),
	.datab(!din_b[189]),
	.datac(!Xd_0__inst_mult_15_177 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_397 ),
	.sharein(Xd_0__inst_mult_15_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_400 ),
	.cout(Xd_0__inst_mult_15_401 ),
	.shareout(Xd_0__inst_mult_15_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_55 (
// Equation(s):
// Xd_0__inst_mult_15_55_sumout  = SUM(( (din_a[190] & din_b[188]) ) + ( Xd_0__inst_mult_6_49  ) + ( Xd_0__inst_mult_6_48  ))
// Xd_0__inst_mult_15_56  = CARRY(( (din_a[190] & din_b[188]) ) + ( Xd_0__inst_mult_6_49  ) + ( Xd_0__inst_mult_6_48  ))
// Xd_0__inst_mult_15_57  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[188]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_48 ),
	.sharein(Xd_0__inst_mult_6_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_55_sumout ),
	.cout(Xd_0__inst_mult_15_56 ),
	.shareout(Xd_0__inst_mult_15_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_115 (
// Equation(s):
// Xd_0__inst_mult_10_372  = SUM(( !Xd_0__inst_mult_10_564  $ (((!din_a[129]) # (!din_b[129]))) ) + ( Xd_0__inst_mult_10_370  ) + ( Xd_0__inst_mult_10_369  ))
// Xd_0__inst_mult_10_373  = CARRY(( !Xd_0__inst_mult_10_564  $ (((!din_a[129]) # (!din_b[129]))) ) + ( Xd_0__inst_mult_10_370  ) + ( Xd_0__inst_mult_10_369  ))
// Xd_0__inst_mult_10_374  = SHARE((din_a[129] & (din_b[129] & Xd_0__inst_mult_10_564 )))

	.dataa(!din_a[129]),
	.datab(!din_b[129]),
	.datac(!Xd_0__inst_mult_10_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_369 ),
	.sharein(Xd_0__inst_mult_10_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_372 ),
	.cout(Xd_0__inst_mult_10_373 ),
	.shareout(Xd_0__inst_mult_10_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_47 (
// Equation(s):
// Xd_0__inst_mult_10_47_sumout  = SUM(( (din_a[130] & din_b[128]) ) + ( Xd_0__inst_mult_11_49  ) + ( Xd_0__inst_mult_11_48  ))
// Xd_0__inst_mult_10_48  = CARRY(( (din_a[130] & din_b[128]) ) + ( Xd_0__inst_mult_11_49  ) + ( Xd_0__inst_mult_11_48  ))
// Xd_0__inst_mult_10_49  = SHARE(GND)

	.dataa(!din_a[130]),
	.datab(!din_b[128]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_48 ),
	.sharein(Xd_0__inst_mult_11_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_47_sumout ),
	.cout(Xd_0__inst_mult_10_48 ),
	.shareout(Xd_0__inst_mult_10_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_119 (
// Equation(s):
// Xd_0__inst_mult_11_376  = SUM(( !Xd_0__inst_mult_11_568  $ (((!din_a[141]) # (!din_b[141]))) ) + ( Xd_0__inst_mult_11_374  ) + ( Xd_0__inst_mult_11_373  ))
// Xd_0__inst_mult_11_377  = CARRY(( !Xd_0__inst_mult_11_568  $ (((!din_a[141]) # (!din_b[141]))) ) + ( Xd_0__inst_mult_11_374  ) + ( Xd_0__inst_mult_11_373  ))
// Xd_0__inst_mult_11_378  = SHARE((din_a[141] & (din_b[141] & Xd_0__inst_mult_11_568 )))

	.dataa(!din_a[141]),
	.datab(!din_b[141]),
	.datac(!Xd_0__inst_mult_11_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_373 ),
	.sharein(Xd_0__inst_mult_11_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_376 ),
	.cout(Xd_0__inst_mult_11_377 ),
	.shareout(Xd_0__inst_mult_11_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_47 (
// Equation(s):
// Xd_0__inst_mult_11_47_sumout  = SUM(( (din_a[142] & din_b[140]) ) + ( Xd_0__inst_mult_8_57  ) + ( Xd_0__inst_mult_8_56  ))
// Xd_0__inst_mult_11_48  = CARRY(( (din_a[142] & din_b[140]) ) + ( Xd_0__inst_mult_8_57  ) + ( Xd_0__inst_mult_8_56  ))
// Xd_0__inst_mult_11_49  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[140]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_56 ),
	.sharein(Xd_0__inst_mult_8_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_47_sumout ),
	.cout(Xd_0__inst_mult_11_48 ),
	.shareout(Xd_0__inst_mult_11_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_119 (
// Equation(s):
// Xd_0__inst_mult_8_376  = SUM(( !Xd_0__inst_mult_8_568  $ (((!din_a[105]) # (!din_b[105]))) ) + ( Xd_0__inst_mult_8_374  ) + ( Xd_0__inst_mult_8_373  ))
// Xd_0__inst_mult_8_377  = CARRY(( !Xd_0__inst_mult_8_568  $ (((!din_a[105]) # (!din_b[105]))) ) + ( Xd_0__inst_mult_8_374  ) + ( Xd_0__inst_mult_8_373  ))
// Xd_0__inst_mult_8_378  = SHARE((din_a[105] & (din_b[105] & Xd_0__inst_mult_8_568 )))

	.dataa(!din_a[105]),
	.datab(!din_b[105]),
	.datac(!Xd_0__inst_mult_8_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_373 ),
	.sharein(Xd_0__inst_mult_8_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_376 ),
	.cout(Xd_0__inst_mult_8_377 ),
	.shareout(Xd_0__inst_mult_8_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_55 (
// Equation(s):
// Xd_0__inst_mult_8_55_sumout  = SUM(( (din_a[106] & din_b[104]) ) + ( Xd_0__inst_mult_9_45  ) + ( Xd_0__inst_mult_9_44  ))
// Xd_0__inst_mult_8_56  = CARRY(( (din_a[106] & din_b[104]) ) + ( Xd_0__inst_mult_9_45  ) + ( Xd_0__inst_mult_9_44  ))
// Xd_0__inst_mult_8_57  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[104]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_44 ),
	.sharein(Xd_0__inst_mult_9_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_55_sumout ),
	.cout(Xd_0__inst_mult_8_56 ),
	.shareout(Xd_0__inst_mult_8_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_115 (
// Equation(s):
// Xd_0__inst_mult_9_372  = SUM(( !Xd_0__inst_mult_9_564  $ (((!din_a[117]) # (!din_b[117]))) ) + ( Xd_0__inst_mult_9_370  ) + ( Xd_0__inst_mult_9_369  ))
// Xd_0__inst_mult_9_373  = CARRY(( !Xd_0__inst_mult_9_564  $ (((!din_a[117]) # (!din_b[117]))) ) + ( Xd_0__inst_mult_9_370  ) + ( Xd_0__inst_mult_9_369  ))
// Xd_0__inst_mult_9_374  = SHARE((din_a[117] & (din_b[117] & Xd_0__inst_mult_9_564 )))

	.dataa(!din_a[117]),
	.datab(!din_b[117]),
	.datac(!Xd_0__inst_mult_9_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_369 ),
	.sharein(Xd_0__inst_mult_9_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_372 ),
	.cout(Xd_0__inst_mult_9_373 ),
	.shareout(Xd_0__inst_mult_9_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_43 (
// Equation(s):
// Xd_0__inst_mult_9_43_sumout  = SUM(( (din_a[118] & din_b[116]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_44  = CARRY(( (din_a[118] & din_b[116]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_45  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[116]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_43_sumout ),
	.cout(Xd_0__inst_mult_9_44 ),
	.shareout(Xd_0__inst_mult_9_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_115 (
// Equation(s):
// Xd_0__inst_mult_6_372  = SUM(( !Xd_0__inst_mult_6_564  $ (((!din_a[81]) # (!din_b[81]))) ) + ( Xd_0__inst_mult_6_370  ) + ( Xd_0__inst_mult_6_369  ))
// Xd_0__inst_mult_6_373  = CARRY(( !Xd_0__inst_mult_6_564  $ (((!din_a[81]) # (!din_b[81]))) ) + ( Xd_0__inst_mult_6_370  ) + ( Xd_0__inst_mult_6_369  ))
// Xd_0__inst_mult_6_374  = SHARE((din_a[81] & (din_b[81] & Xd_0__inst_mult_6_564 )))

	.dataa(!din_a[81]),
	.datab(!din_b[81]),
	.datac(!Xd_0__inst_mult_6_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_369 ),
	.sharein(Xd_0__inst_mult_6_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_372 ),
	.cout(Xd_0__inst_mult_6_373 ),
	.shareout(Xd_0__inst_mult_6_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_51 (
// Equation(s):
// Xd_0__inst_mult_6_51_sumout  = SUM(( (din_a[82] & din_b[80]) ) + ( Xd_0__inst_mult_7_45  ) + ( Xd_0__inst_mult_7_44  ))
// Xd_0__inst_mult_6_52  = CARRY(( (din_a[82] & din_b[80]) ) + ( Xd_0__inst_mult_7_45  ) + ( Xd_0__inst_mult_7_44  ))
// Xd_0__inst_mult_6_53  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_44 ),
	.sharein(Xd_0__inst_mult_7_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_51_sumout ),
	.cout(Xd_0__inst_mult_6_52 ),
	.shareout(Xd_0__inst_mult_6_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_113 (
// Equation(s):
// Xd_0__inst_mult_7_364  = SUM(( !Xd_0__inst_mult_7_564  $ (((!din_a[93]) # (!din_b[93]))) ) + ( Xd_0__inst_mult_7_362  ) + ( Xd_0__inst_mult_7_361  ))
// Xd_0__inst_mult_7_365  = CARRY(( !Xd_0__inst_mult_7_564  $ (((!din_a[93]) # (!din_b[93]))) ) + ( Xd_0__inst_mult_7_362  ) + ( Xd_0__inst_mult_7_361  ))
// Xd_0__inst_mult_7_366  = SHARE((din_a[93] & (din_b[93] & Xd_0__inst_mult_7_564 )))

	.dataa(!din_a[93]),
	.datab(!din_b[93]),
	.datac(!Xd_0__inst_mult_7_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_361 ),
	.sharein(Xd_0__inst_mult_7_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_364 ),
	.cout(Xd_0__inst_mult_7_365 ),
	.shareout(Xd_0__inst_mult_7_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_43 (
// Equation(s):
// Xd_0__inst_mult_7_43_sumout  = SUM(( (din_a[94] & din_b[92]) ) + ( Xd_0__inst_mult_4_49  ) + ( Xd_0__inst_mult_4_48  ))
// Xd_0__inst_mult_7_44  = CARRY(( (din_a[94] & din_b[92]) ) + ( Xd_0__inst_mult_4_49  ) + ( Xd_0__inst_mult_4_48  ))
// Xd_0__inst_mult_7_45  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_48 ),
	.sharein(Xd_0__inst_mult_4_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_43_sumout ),
	.cout(Xd_0__inst_mult_7_44 ),
	.shareout(Xd_0__inst_mult_7_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_125 (
// Equation(s):
// Xd_0__inst_mult_4_400  = SUM(( !Xd_0__inst_mult_4_177  $ (((!din_a[57]) # (!din_b[57]))) ) + ( Xd_0__inst_mult_4_398  ) + ( Xd_0__inst_mult_4_397  ))
// Xd_0__inst_mult_4_401  = CARRY(( !Xd_0__inst_mult_4_177  $ (((!din_a[57]) # (!din_b[57]))) ) + ( Xd_0__inst_mult_4_398  ) + ( Xd_0__inst_mult_4_397  ))
// Xd_0__inst_mult_4_402  = SHARE((din_a[57] & (din_b[57] & Xd_0__inst_mult_4_177 )))

	.dataa(!din_a[57]),
	.datab(!din_b[57]),
	.datac(!Xd_0__inst_mult_4_177 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_397 ),
	.sharein(Xd_0__inst_mult_4_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_400 ),
	.cout(Xd_0__inst_mult_4_401 ),
	.shareout(Xd_0__inst_mult_4_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_47 (
// Equation(s):
// Xd_0__inst_mult_4_47_sumout  = SUM(( (din_a[58] & din_b[56]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_48  = CARRY(( (din_a[58] & din_b[56]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_49  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_47_sumout ),
	.cout(Xd_0__inst_mult_4_48 ),
	.shareout(Xd_0__inst_mult_4_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_113 (
// Equation(s):
// Xd_0__inst_mult_5_364  = SUM(( !Xd_0__inst_mult_5_564  $ (((!din_a[69]) # (!din_b[69]))) ) + ( Xd_0__inst_mult_5_362  ) + ( Xd_0__inst_mult_5_361  ))
// Xd_0__inst_mult_5_365  = CARRY(( !Xd_0__inst_mult_5_564  $ (((!din_a[69]) # (!din_b[69]))) ) + ( Xd_0__inst_mult_5_362  ) + ( Xd_0__inst_mult_5_361  ))
// Xd_0__inst_mult_5_366  = SHARE((din_a[69] & (din_b[69] & Xd_0__inst_mult_5_564 )))

	.dataa(!din_a[69]),
	.datab(!din_b[69]),
	.datac(!Xd_0__inst_mult_5_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_361 ),
	.sharein(Xd_0__inst_mult_5_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_364 ),
	.cout(Xd_0__inst_mult_5_365 ),
	.shareout(Xd_0__inst_mult_5_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_51 (
// Equation(s):
// Xd_0__inst_mult_5_51_sumout  = SUM(( (din_a[70] & din_b[68]) ) + ( Xd_0__inst_mult_8_61  ) + ( Xd_0__inst_mult_8_60  ))
// Xd_0__inst_mult_5_52  = CARRY(( (din_a[70] & din_b[68]) ) + ( Xd_0__inst_mult_8_61  ) + ( Xd_0__inst_mult_8_60  ))
// Xd_0__inst_mult_5_53  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_60 ),
	.sharein(Xd_0__inst_mult_8_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_51_sumout ),
	.cout(Xd_0__inst_mult_5_52 ),
	.shareout(Xd_0__inst_mult_5_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_117 (
// Equation(s):
// Xd_0__inst_mult_2_368  = SUM(( !Xd_0__inst_mult_2_568  $ (((!din_a[33]) # (!din_b[33]))) ) + ( Xd_0__inst_mult_2_366  ) + ( Xd_0__inst_mult_2_365  ))
// Xd_0__inst_mult_2_369  = CARRY(( !Xd_0__inst_mult_2_568  $ (((!din_a[33]) # (!din_b[33]))) ) + ( Xd_0__inst_mult_2_366  ) + ( Xd_0__inst_mult_2_365  ))
// Xd_0__inst_mult_2_370  = SHARE((din_a[33] & (din_b[33] & Xd_0__inst_mult_2_568 )))

	.dataa(!din_a[33]),
	.datab(!din_b[33]),
	.datac(!Xd_0__inst_mult_2_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_365 ),
	.sharein(Xd_0__inst_mult_2_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_368 ),
	.cout(Xd_0__inst_mult_2_369 ),
	.shareout(Xd_0__inst_mult_2_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_51 (
// Equation(s):
// Xd_0__inst_mult_2_51_sumout  = SUM(( (din_a[34] & din_b[32]) ) + ( Xd_0__inst_mult_3_57  ) + ( Xd_0__inst_mult_3_56  ))
// Xd_0__inst_mult_2_52  = CARRY(( (din_a[34] & din_b[32]) ) + ( Xd_0__inst_mult_3_57  ) + ( Xd_0__inst_mult_3_56  ))
// Xd_0__inst_mult_2_53  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_56 ),
	.sharein(Xd_0__inst_mult_3_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_51_sumout ),
	.cout(Xd_0__inst_mult_2_52 ),
	.shareout(Xd_0__inst_mult_2_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_113 (
// Equation(s):
// Xd_0__inst_mult_3_364  = SUM(( !Xd_0__inst_mult_3_564  $ (((!din_a[45]) # (!din_b[45]))) ) + ( Xd_0__inst_mult_3_362  ) + ( Xd_0__inst_mult_3_361  ))
// Xd_0__inst_mult_3_365  = CARRY(( !Xd_0__inst_mult_3_564  $ (((!din_a[45]) # (!din_b[45]))) ) + ( Xd_0__inst_mult_3_362  ) + ( Xd_0__inst_mult_3_361  ))
// Xd_0__inst_mult_3_366  = SHARE((din_a[45] & (din_b[45] & Xd_0__inst_mult_3_564 )))

	.dataa(!din_a[45]),
	.datab(!din_b[45]),
	.datac(!Xd_0__inst_mult_3_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_361 ),
	.sharein(Xd_0__inst_mult_3_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_364 ),
	.cout(Xd_0__inst_mult_3_365 ),
	.shareout(Xd_0__inst_mult_3_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_55 (
// Equation(s):
// Xd_0__inst_mult_3_55_sumout  = SUM(( (din_a[46] & din_b[44]) ) + ( Xd_0__inst_mult_0_49  ) + ( Xd_0__inst_mult_0_48  ))
// Xd_0__inst_mult_3_56  = CARRY(( (din_a[46] & din_b[44]) ) + ( Xd_0__inst_mult_0_49  ) + ( Xd_0__inst_mult_0_48  ))
// Xd_0__inst_mult_3_57  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_48 ),
	.sharein(Xd_0__inst_mult_0_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_55_sumout ),
	.cout(Xd_0__inst_mult_3_56 ),
	.shareout(Xd_0__inst_mult_3_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_118 (
// Equation(s):
// Xd_0__inst_mult_0_372  = SUM(( !Xd_0__inst_mult_0_568  $ (((!din_a[9]) # (!din_b[9]))) ) + ( Xd_0__inst_mult_0_370  ) + ( Xd_0__inst_mult_0_369  ))
// Xd_0__inst_mult_0_373  = CARRY(( !Xd_0__inst_mult_0_568  $ (((!din_a[9]) # (!din_b[9]))) ) + ( Xd_0__inst_mult_0_370  ) + ( Xd_0__inst_mult_0_369  ))
// Xd_0__inst_mult_0_374  = SHARE((din_a[9] & (din_b[9] & Xd_0__inst_mult_0_568 )))

	.dataa(!din_a[9]),
	.datab(!din_b[9]),
	.datac(!Xd_0__inst_mult_0_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_369 ),
	.sharein(Xd_0__inst_mult_0_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_372 ),
	.cout(Xd_0__inst_mult_0_373 ),
	.shareout(Xd_0__inst_mult_0_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_47 (
// Equation(s):
// Xd_0__inst_mult_0_47_sumout  = SUM(( (din_a[10] & din_b[8]) ) + ( Xd_0__inst_mult_1_53  ) + ( Xd_0__inst_mult_1_52  ))
// Xd_0__inst_mult_0_48  = CARRY(( (din_a[10] & din_b[8]) ) + ( Xd_0__inst_mult_1_53  ) + ( Xd_0__inst_mult_1_52  ))
// Xd_0__inst_mult_0_49  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_52 ),
	.sharein(Xd_0__inst_mult_1_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_47_sumout ),
	.cout(Xd_0__inst_mult_0_48 ),
	.shareout(Xd_0__inst_mult_0_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_118 (
// Equation(s):
// Xd_0__inst_mult_1_372  = SUM(( !Xd_0__inst_mult_1_572  $ (((!din_a[21]) # (!din_b[21]))) ) + ( Xd_0__inst_mult_1_370  ) + ( Xd_0__inst_mult_1_369  ))
// Xd_0__inst_mult_1_373  = CARRY(( !Xd_0__inst_mult_1_572  $ (((!din_a[21]) # (!din_b[21]))) ) + ( Xd_0__inst_mult_1_370  ) + ( Xd_0__inst_mult_1_369  ))
// Xd_0__inst_mult_1_374  = SHARE((din_a[21] & (din_b[21] & Xd_0__inst_mult_1_572 )))

	.dataa(!din_a[21]),
	.datab(!din_b[21]),
	.datac(!Xd_0__inst_mult_1_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_369 ),
	.sharein(Xd_0__inst_mult_1_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_372 ),
	.cout(Xd_0__inst_mult_1_373 ),
	.shareout(Xd_0__inst_mult_1_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_51 (
// Equation(s):
// Xd_0__inst_mult_1_51_sumout  = SUM(( (din_a[22] & din_b[20]) ) + ( Xd_0__inst_mult_14_65  ) + ( Xd_0__inst_mult_14_64  ))
// Xd_0__inst_mult_1_52  = CARRY(( (din_a[22] & din_b[20]) ) + ( Xd_0__inst_mult_14_65  ) + ( Xd_0__inst_mult_14_64  ))
// Xd_0__inst_mult_1_53  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_64 ),
	.sharein(Xd_0__inst_mult_14_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_51_sumout ),
	.cout(Xd_0__inst_mult_1_52 ),
	.shareout(Xd_0__inst_mult_1_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_122 (
// Equation(s):
// Xd_0__inst_mult_12_400  = SUM(( !Xd_0__inst_mult_12_169  $ (((!din_a[153]) # (!din_b[154]))) ) + ( Xd_0__inst_mult_12_398  ) + ( Xd_0__inst_mult_12_397  ))
// Xd_0__inst_mult_12_401  = CARRY(( !Xd_0__inst_mult_12_169  $ (((!din_a[153]) # (!din_b[154]))) ) + ( Xd_0__inst_mult_12_398  ) + ( Xd_0__inst_mult_12_397  ))
// Xd_0__inst_mult_12_402  = SHARE((din_a[153] & (din_b[154] & Xd_0__inst_mult_12_169 )))

	.dataa(!din_a[153]),
	.datab(!din_b[154]),
	.datac(!Xd_0__inst_mult_12_169 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_397 ),
	.sharein(Xd_0__inst_mult_12_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_400 ),
	.cout(Xd_0__inst_mult_12_401 ),
	.shareout(Xd_0__inst_mult_12_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_59 (
// Equation(s):
// Xd_0__inst_mult_12_59_sumout  = SUM(( (din_a[154] & din_b[153]) ) + ( Xd_0__inst_mult_13_57  ) + ( Xd_0__inst_mult_13_56  ))
// Xd_0__inst_mult_12_60  = CARRY(( (din_a[154] & din_b[153]) ) + ( Xd_0__inst_mult_13_57  ) + ( Xd_0__inst_mult_13_56  ))
// Xd_0__inst_mult_12_61  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[153]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_56 ),
	.sharein(Xd_0__inst_mult_13_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_59_sumout ),
	.cout(Xd_0__inst_mult_12_60 ),
	.shareout(Xd_0__inst_mult_12_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_120 (
// Equation(s):
// Xd_0__inst_mult_13_380  = SUM(( !Xd_0__inst_mult_13_572  $ (((!din_a[165]) # (!din_b[166]))) ) + ( Xd_0__inst_mult_13_378  ) + ( Xd_0__inst_mult_13_377  ))
// Xd_0__inst_mult_13_381  = CARRY(( !Xd_0__inst_mult_13_572  $ (((!din_a[165]) # (!din_b[166]))) ) + ( Xd_0__inst_mult_13_378  ) + ( Xd_0__inst_mult_13_377  ))
// Xd_0__inst_mult_13_382  = SHARE((din_a[165] & (din_b[166] & Xd_0__inst_mult_13_572 )))

	.dataa(!din_a[165]),
	.datab(!din_b[166]),
	.datac(!Xd_0__inst_mult_13_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_377 ),
	.sharein(Xd_0__inst_mult_13_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_380 ),
	.cout(Xd_0__inst_mult_13_381 ),
	.shareout(Xd_0__inst_mult_13_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_55 (
// Equation(s):
// Xd_0__inst_mult_13_55_sumout  = SUM(( (din_a[166] & din_b[165]) ) + ( Xd_0__inst_mult_10_53  ) + ( Xd_0__inst_mult_10_52  ))
// Xd_0__inst_mult_13_56  = CARRY(( (din_a[166] & din_b[165]) ) + ( Xd_0__inst_mult_10_53  ) + ( Xd_0__inst_mult_10_52  ))
// Xd_0__inst_mult_13_57  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[165]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_52 ),
	.sharein(Xd_0__inst_mult_10_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_55_sumout ),
	.cout(Xd_0__inst_mult_13_56 ),
	.shareout(Xd_0__inst_mult_13_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_124 (
// Equation(s):
// Xd_0__inst_mult_14_396  = SUM(( !Xd_0__inst_mult_14_576  $ (((!din_a[177]) # (!din_b[178]))) ) + ( Xd_0__inst_mult_14_394  ) + ( Xd_0__inst_mult_14_393  ))
// Xd_0__inst_mult_14_397  = CARRY(( !Xd_0__inst_mult_14_576  $ (((!din_a[177]) # (!din_b[178]))) ) + ( Xd_0__inst_mult_14_394  ) + ( Xd_0__inst_mult_14_393  ))
// Xd_0__inst_mult_14_398  = SHARE((din_a[177] & (din_b[178] & Xd_0__inst_mult_14_576 )))

	.dataa(!din_a[177]),
	.datab(!din_b[178]),
	.datac(!Xd_0__inst_mult_14_576 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_393 ),
	.sharein(Xd_0__inst_mult_14_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_396 ),
	.cout(Xd_0__inst_mult_14_397 ),
	.shareout(Xd_0__inst_mult_14_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_63 (
// Equation(s):
// Xd_0__inst_mult_14_63_sumout  = SUM(( (din_a[178] & din_b[177]) ) + ( Xd_0__inst_mult_15_61  ) + ( Xd_0__inst_mult_15_60  ))
// Xd_0__inst_mult_14_64  = CARRY(( (din_a[178] & din_b[177]) ) + ( Xd_0__inst_mult_15_61  ) + ( Xd_0__inst_mult_15_60  ))
// Xd_0__inst_mult_14_65  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[177]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_60 ),
	.sharein(Xd_0__inst_mult_15_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_63_sumout ),
	.cout(Xd_0__inst_mult_14_64 ),
	.shareout(Xd_0__inst_mult_14_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_126 (
// Equation(s):
// Xd_0__inst_mult_15_404  = SUM(( !Xd_0__inst_mult_15_173  $ (((!din_a[189]) # (!din_b[190]))) ) + ( Xd_0__inst_mult_15_402  ) + ( Xd_0__inst_mult_15_401  ))
// Xd_0__inst_mult_15_405  = CARRY(( !Xd_0__inst_mult_15_173  $ (((!din_a[189]) # (!din_b[190]))) ) + ( Xd_0__inst_mult_15_402  ) + ( Xd_0__inst_mult_15_401  ))
// Xd_0__inst_mult_15_406  = SHARE((din_a[189] & (din_b[190] & Xd_0__inst_mult_15_173 )))

	.dataa(!din_a[189]),
	.datab(!din_b[190]),
	.datac(!Xd_0__inst_mult_15_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_401 ),
	.sharein(Xd_0__inst_mult_15_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_404 ),
	.cout(Xd_0__inst_mult_15_405 ),
	.shareout(Xd_0__inst_mult_15_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_59 (
// Equation(s):
// Xd_0__inst_mult_15_59_sumout  = SUM(( (din_a[190] & din_b[189]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_60  = CARRY(( (din_a[190] & din_b[189]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_61  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[189]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_15_59_sumout ),
	.cout(Xd_0__inst_mult_15_60 ),
	.shareout(Xd_0__inst_mult_15_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_116 (
// Equation(s):
// Xd_0__inst_mult_10_376  = SUM(( !Xd_0__inst_mult_10_568  $ (((!din_a[129]) # (!din_b[130]))) ) + ( Xd_0__inst_mult_10_374  ) + ( Xd_0__inst_mult_10_373  ))
// Xd_0__inst_mult_10_377  = CARRY(( !Xd_0__inst_mult_10_568  $ (((!din_a[129]) # (!din_b[130]))) ) + ( Xd_0__inst_mult_10_374  ) + ( Xd_0__inst_mult_10_373  ))
// Xd_0__inst_mult_10_378  = SHARE((din_a[129] & (din_b[130] & Xd_0__inst_mult_10_568 )))

	.dataa(!din_a[129]),
	.datab(!din_b[130]),
	.datac(!Xd_0__inst_mult_10_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_373 ),
	.sharein(Xd_0__inst_mult_10_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_376 ),
	.cout(Xd_0__inst_mult_10_377 ),
	.shareout(Xd_0__inst_mult_10_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_51 (
// Equation(s):
// Xd_0__inst_mult_10_51_sumout  = SUM(( (din_a[130] & din_b[129]) ) + ( Xd_0__inst_mult_5_53  ) + ( Xd_0__inst_mult_5_52  ))
// Xd_0__inst_mult_10_52  = CARRY(( (din_a[130] & din_b[129]) ) + ( Xd_0__inst_mult_5_53  ) + ( Xd_0__inst_mult_5_52  ))
// Xd_0__inst_mult_10_53  = SHARE(GND)

	.dataa(!din_a[130]),
	.datab(!din_b[129]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_52 ),
	.sharein(Xd_0__inst_mult_5_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_51_sumout ),
	.cout(Xd_0__inst_mult_10_52 ),
	.shareout(Xd_0__inst_mult_10_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_120 (
// Equation(s):
// Xd_0__inst_mult_11_380  = SUM(( !Xd_0__inst_mult_11_572  $ (((!din_a[141]) # (!din_b[142]))) ) + ( Xd_0__inst_mult_11_378  ) + ( Xd_0__inst_mult_11_377  ))
// Xd_0__inst_mult_11_381  = CARRY(( !Xd_0__inst_mult_11_572  $ (((!din_a[141]) # (!din_b[142]))) ) + ( Xd_0__inst_mult_11_378  ) + ( Xd_0__inst_mult_11_377  ))
// Xd_0__inst_mult_11_382  = SHARE((din_a[141] & (din_b[142] & Xd_0__inst_mult_11_572 )))

	.dataa(!din_a[141]),
	.datab(!din_b[142]),
	.datac(!Xd_0__inst_mult_11_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_377 ),
	.sharein(Xd_0__inst_mult_11_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_380 ),
	.cout(Xd_0__inst_mult_11_381 ),
	.shareout(Xd_0__inst_mult_11_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_51 (
// Equation(s):
// Xd_0__inst_mult_11_51_sumout  = SUM(( (din_a[142] & din_b[141]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_52  = CARRY(( (din_a[142] & din_b[141]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_53  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[141]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_51_sumout ),
	.cout(Xd_0__inst_mult_11_52 ),
	.shareout(Xd_0__inst_mult_11_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_120 (
// Equation(s):
// Xd_0__inst_mult_8_380  = SUM(( !Xd_0__inst_mult_8_572  $ (((!din_a[105]) # (!din_b[106]))) ) + ( Xd_0__inst_mult_8_378  ) + ( Xd_0__inst_mult_8_377  ))
// Xd_0__inst_mult_8_381  = CARRY(( !Xd_0__inst_mult_8_572  $ (((!din_a[105]) # (!din_b[106]))) ) + ( Xd_0__inst_mult_8_378  ) + ( Xd_0__inst_mult_8_377  ))
// Xd_0__inst_mult_8_382  = SHARE((din_a[105] & (din_b[106] & Xd_0__inst_mult_8_572 )))

	.dataa(!din_a[105]),
	.datab(!din_b[106]),
	.datac(!Xd_0__inst_mult_8_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_377 ),
	.sharein(Xd_0__inst_mult_8_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_380 ),
	.cout(Xd_0__inst_mult_8_381 ),
	.shareout(Xd_0__inst_mult_8_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_59 (
// Equation(s):
// Xd_0__inst_mult_8_59_sumout  = SUM(( (din_a[106] & din_b[105]) ) + ( Xd_0__inst_mult_9_49  ) + ( Xd_0__inst_mult_9_48  ))
// Xd_0__inst_mult_8_60  = CARRY(( (din_a[106] & din_b[105]) ) + ( Xd_0__inst_mult_9_49  ) + ( Xd_0__inst_mult_9_48  ))
// Xd_0__inst_mult_8_61  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[105]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_48 ),
	.sharein(Xd_0__inst_mult_9_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_59_sumout ),
	.cout(Xd_0__inst_mult_8_60 ),
	.shareout(Xd_0__inst_mult_8_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_116 (
// Equation(s):
// Xd_0__inst_mult_9_376  = SUM(( !Xd_0__inst_mult_9_568  $ (((!din_a[117]) # (!din_b[118]))) ) + ( Xd_0__inst_mult_9_374  ) + ( Xd_0__inst_mult_9_373  ))
// Xd_0__inst_mult_9_377  = CARRY(( !Xd_0__inst_mult_9_568  $ (((!din_a[117]) # (!din_b[118]))) ) + ( Xd_0__inst_mult_9_374  ) + ( Xd_0__inst_mult_9_373  ))
// Xd_0__inst_mult_9_378  = SHARE((din_a[117] & (din_b[118] & Xd_0__inst_mult_9_568 )))

	.dataa(!din_a[117]),
	.datab(!din_b[118]),
	.datac(!Xd_0__inst_mult_9_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_373 ),
	.sharein(Xd_0__inst_mult_9_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_376 ),
	.cout(Xd_0__inst_mult_9_377 ),
	.shareout(Xd_0__inst_mult_9_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_47 (
// Equation(s):
// Xd_0__inst_mult_9_47_sumout  = SUM(( (din_a[118] & din_b[117]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_48  = CARRY(( (din_a[118] & din_b[117]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_49  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[117]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_47_sumout ),
	.cout(Xd_0__inst_mult_9_48 ),
	.shareout(Xd_0__inst_mult_9_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_116 (
// Equation(s):
// Xd_0__inst_mult_6_376  = SUM(( !Xd_0__inst_mult_6_568  $ (((!din_a[81]) # (!din_b[82]))) ) + ( Xd_0__inst_mult_6_374  ) + ( Xd_0__inst_mult_6_373  ))
// Xd_0__inst_mult_6_377  = CARRY(( !Xd_0__inst_mult_6_568  $ (((!din_a[81]) # (!din_b[82]))) ) + ( Xd_0__inst_mult_6_374  ) + ( Xd_0__inst_mult_6_373  ))
// Xd_0__inst_mult_6_378  = SHARE((din_a[81] & (din_b[82] & Xd_0__inst_mult_6_568 )))

	.dataa(!din_a[81]),
	.datab(!din_b[82]),
	.datac(!Xd_0__inst_mult_6_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_373 ),
	.sharein(Xd_0__inst_mult_6_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_376 ),
	.cout(Xd_0__inst_mult_6_377 ),
	.shareout(Xd_0__inst_mult_6_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_55 (
// Equation(s):
// Xd_0__inst_mult_6_55_sumout  = SUM(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_7_49  ) + ( Xd_0__inst_mult_7_48  ))
// Xd_0__inst_mult_6_56  = CARRY(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_7_49  ) + ( Xd_0__inst_mult_7_48  ))
// Xd_0__inst_mult_6_57  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[81]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_48 ),
	.sharein(Xd_0__inst_mult_7_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_55_sumout ),
	.cout(Xd_0__inst_mult_6_56 ),
	.shareout(Xd_0__inst_mult_6_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_114 (
// Equation(s):
// Xd_0__inst_mult_7_368  = SUM(( !Xd_0__inst_mult_7_568  $ (((!din_a[93]) # (!din_b[94]))) ) + ( Xd_0__inst_mult_7_366  ) + ( Xd_0__inst_mult_7_365  ))
// Xd_0__inst_mult_7_369  = CARRY(( !Xd_0__inst_mult_7_568  $ (((!din_a[93]) # (!din_b[94]))) ) + ( Xd_0__inst_mult_7_366  ) + ( Xd_0__inst_mult_7_365  ))
// Xd_0__inst_mult_7_370  = SHARE((din_a[93] & (din_b[94] & Xd_0__inst_mult_7_568 )))

	.dataa(!din_a[93]),
	.datab(!din_b[94]),
	.datac(!Xd_0__inst_mult_7_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_365 ),
	.sharein(Xd_0__inst_mult_7_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_368 ),
	.cout(Xd_0__inst_mult_7_369 ),
	.shareout(Xd_0__inst_mult_7_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_47 (
// Equation(s):
// Xd_0__inst_mult_7_47_sumout  = SUM(( (din_a[94] & din_b[93]) ) + ( Xd_0__inst_mult_4_53  ) + ( Xd_0__inst_mult_4_52  ))
// Xd_0__inst_mult_7_48  = CARRY(( (din_a[94] & din_b[93]) ) + ( Xd_0__inst_mult_4_53  ) + ( Xd_0__inst_mult_4_52  ))
// Xd_0__inst_mult_7_49  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_52 ),
	.sharein(Xd_0__inst_mult_4_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_47_sumout ),
	.cout(Xd_0__inst_mult_7_48 ),
	.shareout(Xd_0__inst_mult_7_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_126 (
// Equation(s):
// Xd_0__inst_mult_4_404  = SUM(( !Xd_0__inst_mult_4_173  $ (((!din_a[57]) # (!din_b[58]))) ) + ( Xd_0__inst_mult_4_402  ) + ( Xd_0__inst_mult_4_401  ))
// Xd_0__inst_mult_4_405  = CARRY(( !Xd_0__inst_mult_4_173  $ (((!din_a[57]) # (!din_b[58]))) ) + ( Xd_0__inst_mult_4_402  ) + ( Xd_0__inst_mult_4_401  ))
// Xd_0__inst_mult_4_406  = SHARE((din_a[57] & (din_b[58] & Xd_0__inst_mult_4_173 )))

	.dataa(!din_a[57]),
	.datab(!din_b[58]),
	.datac(!Xd_0__inst_mult_4_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_401 ),
	.sharein(Xd_0__inst_mult_4_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_404 ),
	.cout(Xd_0__inst_mult_4_405 ),
	.shareout(Xd_0__inst_mult_4_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_51 (
// Equation(s):
// Xd_0__inst_mult_4_51_sumout  = SUM(( (din_a[58] & din_b[57]) ) + ( Xd_0__inst_mult_5_57  ) + ( Xd_0__inst_mult_5_56  ))
// Xd_0__inst_mult_4_52  = CARRY(( (din_a[58] & din_b[57]) ) + ( Xd_0__inst_mult_5_57  ) + ( Xd_0__inst_mult_5_56  ))
// Xd_0__inst_mult_4_53  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[57]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_56 ),
	.sharein(Xd_0__inst_mult_5_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_51_sumout ),
	.cout(Xd_0__inst_mult_4_52 ),
	.shareout(Xd_0__inst_mult_4_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_114 (
// Equation(s):
// Xd_0__inst_mult_5_368  = SUM(( !Xd_0__inst_mult_5_568  $ (((!din_a[69]) # (!din_b[70]))) ) + ( Xd_0__inst_mult_5_366  ) + ( Xd_0__inst_mult_5_365  ))
// Xd_0__inst_mult_5_369  = CARRY(( !Xd_0__inst_mult_5_568  $ (((!din_a[69]) # (!din_b[70]))) ) + ( Xd_0__inst_mult_5_366  ) + ( Xd_0__inst_mult_5_365  ))
// Xd_0__inst_mult_5_370  = SHARE((din_a[69] & (din_b[70] & Xd_0__inst_mult_5_568 )))

	.dataa(!din_a[69]),
	.datab(!din_b[70]),
	.datac(!Xd_0__inst_mult_5_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_365 ),
	.sharein(Xd_0__inst_mult_5_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_368 ),
	.cout(Xd_0__inst_mult_5_369 ),
	.shareout(Xd_0__inst_mult_5_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_55 (
// Equation(s):
// Xd_0__inst_mult_5_55_sumout  = SUM(( (din_a[70] & din_b[69]) ) + ( Xd_0__inst_mult_2_57  ) + ( Xd_0__inst_mult_2_56  ))
// Xd_0__inst_mult_5_56  = CARRY(( (din_a[70] & din_b[69]) ) + ( Xd_0__inst_mult_2_57  ) + ( Xd_0__inst_mult_2_56  ))
// Xd_0__inst_mult_5_57  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_56 ),
	.sharein(Xd_0__inst_mult_2_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_55_sumout ),
	.cout(Xd_0__inst_mult_5_56 ),
	.shareout(Xd_0__inst_mult_5_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_118 (
// Equation(s):
// Xd_0__inst_mult_2_372  = SUM(( !Xd_0__inst_mult_2_572  $ (((!din_a[33]) # (!din_b[34]))) ) + ( Xd_0__inst_mult_2_370  ) + ( Xd_0__inst_mult_2_369  ))
// Xd_0__inst_mult_2_373  = CARRY(( !Xd_0__inst_mult_2_572  $ (((!din_a[33]) # (!din_b[34]))) ) + ( Xd_0__inst_mult_2_370  ) + ( Xd_0__inst_mult_2_369  ))
// Xd_0__inst_mult_2_374  = SHARE((din_a[33] & (din_b[34] & Xd_0__inst_mult_2_572 )))

	.dataa(!din_a[33]),
	.datab(!din_b[34]),
	.datac(!Xd_0__inst_mult_2_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_369 ),
	.sharein(Xd_0__inst_mult_2_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_372 ),
	.cout(Xd_0__inst_mult_2_373 ),
	.shareout(Xd_0__inst_mult_2_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_55 (
// Equation(s):
// Xd_0__inst_mult_2_55_sumout  = SUM(( (din_a[34] & din_b[33]) ) + ( Xd_0__inst_mult_3_61  ) + ( Xd_0__inst_mult_3_60  ))
// Xd_0__inst_mult_2_56  = CARRY(( (din_a[34] & din_b[33]) ) + ( Xd_0__inst_mult_3_61  ) + ( Xd_0__inst_mult_3_60  ))
// Xd_0__inst_mult_2_57  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[33]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_60 ),
	.sharein(Xd_0__inst_mult_3_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_55_sumout ),
	.cout(Xd_0__inst_mult_2_56 ),
	.shareout(Xd_0__inst_mult_2_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_114 (
// Equation(s):
// Xd_0__inst_mult_3_368  = SUM(( !Xd_0__inst_mult_3_568  $ (((!din_a[45]) # (!din_b[46]))) ) + ( Xd_0__inst_mult_3_366  ) + ( Xd_0__inst_mult_3_365  ))
// Xd_0__inst_mult_3_369  = CARRY(( !Xd_0__inst_mult_3_568  $ (((!din_a[45]) # (!din_b[46]))) ) + ( Xd_0__inst_mult_3_366  ) + ( Xd_0__inst_mult_3_365  ))
// Xd_0__inst_mult_3_370  = SHARE((din_a[45] & (din_b[46] & Xd_0__inst_mult_3_568 )))

	.dataa(!din_a[45]),
	.datab(!din_b[46]),
	.datac(!Xd_0__inst_mult_3_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_365 ),
	.sharein(Xd_0__inst_mult_3_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_368 ),
	.cout(Xd_0__inst_mult_3_369 ),
	.shareout(Xd_0__inst_mult_3_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_59 (
// Equation(s):
// Xd_0__inst_mult_3_59_sumout  = SUM(( (din_a[46] & din_b[45]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_60  = CARRY(( (din_a[46] & din_b[45]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_61  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[45]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_59_sumout ),
	.cout(Xd_0__inst_mult_3_60 ),
	.shareout(Xd_0__inst_mult_3_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_119 (
// Equation(s):
// Xd_0__inst_mult_0_376  = SUM(( !Xd_0__inst_mult_0_572  $ (((!din_a[9]) # (!din_b[10]))) ) + ( Xd_0__inst_mult_0_374  ) + ( Xd_0__inst_mult_0_373  ))
// Xd_0__inst_mult_0_377  = CARRY(( !Xd_0__inst_mult_0_572  $ (((!din_a[9]) # (!din_b[10]))) ) + ( Xd_0__inst_mult_0_374  ) + ( Xd_0__inst_mult_0_373  ))
// Xd_0__inst_mult_0_378  = SHARE((din_a[9] & (din_b[10] & Xd_0__inst_mult_0_572 )))

	.dataa(!din_a[9]),
	.datab(!din_b[10]),
	.datac(!Xd_0__inst_mult_0_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_373 ),
	.sharein(Xd_0__inst_mult_0_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_376 ),
	.cout(Xd_0__inst_mult_0_377 ),
	.shareout(Xd_0__inst_mult_0_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_51 (
// Equation(s):
// Xd_0__inst_mult_0_51_sumout  = SUM(( (din_a[10] & din_b[9]) ) + ( Xd_0__inst_mult_15_57  ) + ( Xd_0__inst_mult_15_56  ))
// Xd_0__inst_mult_0_52  = CARRY(( (din_a[10] & din_b[9]) ) + ( Xd_0__inst_mult_15_57  ) + ( Xd_0__inst_mult_15_56  ))
// Xd_0__inst_mult_0_53  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[9]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_56 ),
	.sharein(Xd_0__inst_mult_15_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_51_sumout ),
	.cout(Xd_0__inst_mult_0_52 ),
	.shareout(Xd_0__inst_mult_0_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_119 (
// Equation(s):
// Xd_0__inst_mult_1_376  = SUM(( !Xd_0__inst_mult_1_576  $ (((!din_a[21]) # (!din_b[22]))) ) + ( Xd_0__inst_mult_1_374  ) + ( Xd_0__inst_mult_1_373  ))
// Xd_0__inst_mult_1_377  = CARRY(( !Xd_0__inst_mult_1_576  $ (((!din_a[21]) # (!din_b[22]))) ) + ( Xd_0__inst_mult_1_374  ) + ( Xd_0__inst_mult_1_373  ))
// Xd_0__inst_mult_1_378  = SHARE((din_a[21] & (din_b[22] & Xd_0__inst_mult_1_576 )))

	.dataa(!din_a[21]),
	.datab(!din_b[22]),
	.datac(!Xd_0__inst_mult_1_576 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_373 ),
	.sharein(Xd_0__inst_mult_1_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_376 ),
	.cout(Xd_0__inst_mult_1_377 ),
	.shareout(Xd_0__inst_mult_1_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_55 (
// Equation(s):
// Xd_0__inst_mult_1_55_sumout  = SUM(( (din_a[22] & din_b[21]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_56  = CARRY(( (din_a[22] & din_b[21]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_57  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[21]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_55_sumout ),
	.cout(Xd_0__inst_mult_1_56 ),
	.shareout(Xd_0__inst_mult_1_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_123 (
// Equation(s):
// Xd_0__inst_mult_12_404  = SUM(( GND ) + ( Xd_0__inst_mult_12_402  ) + ( Xd_0__inst_mult_12_401  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_401 ),
	.sharein(Xd_0__inst_mult_12_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_404 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_121 (
// Equation(s):
// Xd_0__inst_mult_13_384  = SUM(( GND ) + ( Xd_0__inst_mult_13_382  ) + ( Xd_0__inst_mult_13_381  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_381 ),
	.sharein(Xd_0__inst_mult_13_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_384 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_59 (
// Equation(s):
// Xd_0__inst_mult_13_59_sumout  = SUM(( (din_a[166] & din_b[166]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_60  = CARRY(( (din_a[166] & din_b[166]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_61  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_13_59_sumout ),
	.cout(Xd_0__inst_mult_13_60 ),
	.shareout(Xd_0__inst_mult_13_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_125 (
// Equation(s):
// Xd_0__inst_mult_14_400  = SUM(( GND ) + ( Xd_0__inst_mult_14_398  ) + ( Xd_0__inst_mult_14_397  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_397 ),
	.sharein(Xd_0__inst_mult_14_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_400 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_127 (
// Equation(s):
// Xd_0__inst_mult_15_408  = SUM(( GND ) + ( Xd_0__inst_mult_15_406  ) + ( Xd_0__inst_mult_15_405  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_405 ),
	.sharein(Xd_0__inst_mult_15_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_408 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_117 (
// Equation(s):
// Xd_0__inst_mult_10_380  = SUM(( GND ) + ( Xd_0__inst_mult_10_378  ) + ( Xd_0__inst_mult_10_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_377 ),
	.sharein(Xd_0__inst_mult_10_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_55 (
// Equation(s):
// Xd_0__inst_mult_10_55_sumout  = SUM(( (din_a[130] & din_b[130]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_56  = CARRY(( (din_a[130] & din_b[130]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_57  = SHARE(GND)

	.dataa(!din_a[130]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_10_55_sumout ),
	.cout(Xd_0__inst_mult_10_56 ),
	.shareout(Xd_0__inst_mult_10_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_121 (
// Equation(s):
// Xd_0__inst_mult_11_384  = SUM(( GND ) + ( Xd_0__inst_mult_11_382  ) + ( Xd_0__inst_mult_11_381  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_381 ),
	.sharein(Xd_0__inst_mult_11_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_384 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_121 (
// Equation(s):
// Xd_0__inst_mult_8_384  = SUM(( GND ) + ( Xd_0__inst_mult_8_382  ) + ( Xd_0__inst_mult_8_381  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_381 ),
	.sharein(Xd_0__inst_mult_8_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_384 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_117 (
// Equation(s):
// Xd_0__inst_mult_9_380  = SUM(( GND ) + ( Xd_0__inst_mult_9_378  ) + ( Xd_0__inst_mult_9_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_377 ),
	.sharein(Xd_0__inst_mult_9_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_51 (
// Equation(s):
// Xd_0__inst_mult_9_51_sumout  = SUM(( (din_a[118] & din_b[118]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_52  = CARRY(( (din_a[118] & din_b[118]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_53  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_51_sumout ),
	.cout(Xd_0__inst_mult_9_52 ),
	.shareout(Xd_0__inst_mult_9_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_117 (
// Equation(s):
// Xd_0__inst_mult_6_380  = SUM(( GND ) + ( Xd_0__inst_mult_6_378  ) + ( Xd_0__inst_mult_6_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_377 ),
	.sharein(Xd_0__inst_mult_6_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_115 (
// Equation(s):
// Xd_0__inst_mult_7_372  = SUM(( GND ) + ( Xd_0__inst_mult_7_370  ) + ( Xd_0__inst_mult_7_369  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_369 ),
	.sharein(Xd_0__inst_mult_7_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_372 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_51 (
// Equation(s):
// Xd_0__inst_mult_7_51_sumout  = SUM(( (din_a[94] & din_b[94]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_52  = CARRY(( (din_a[94] & din_b[94]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_53  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_51_sumout ),
	.cout(Xd_0__inst_mult_7_52 ),
	.shareout(Xd_0__inst_mult_7_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_127 (
// Equation(s):
// Xd_0__inst_mult_4_408  = SUM(( GND ) + ( Xd_0__inst_mult_4_406  ) + ( Xd_0__inst_mult_4_405  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_405 ),
	.sharein(Xd_0__inst_mult_4_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_408 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_115 (
// Equation(s):
// Xd_0__inst_mult_5_372  = SUM(( GND ) + ( Xd_0__inst_mult_5_370  ) + ( Xd_0__inst_mult_5_369  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_369 ),
	.sharein(Xd_0__inst_mult_5_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_372 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_119 (
// Equation(s):
// Xd_0__inst_mult_2_376  = SUM(( GND ) + ( Xd_0__inst_mult_2_374  ) + ( Xd_0__inst_mult_2_373  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_373 ),
	.sharein(Xd_0__inst_mult_2_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_376 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_115 (
// Equation(s):
// Xd_0__inst_mult_3_372  = SUM(( GND ) + ( Xd_0__inst_mult_3_370  ) + ( Xd_0__inst_mult_3_369  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_369 ),
	.sharein(Xd_0__inst_mult_3_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_372 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_120 (
// Equation(s):
// Xd_0__inst_mult_0_380  = SUM(( GND ) + ( Xd_0__inst_mult_0_378  ) + ( Xd_0__inst_mult_0_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_377 ),
	.sharein(Xd_0__inst_mult_0_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_55 (
// Equation(s):
// Xd_0__inst_mult_0_55_sumout  = SUM(( (din_a[10] & din_b[10]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_56  = CARRY(( (din_a[10] & din_b[10]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_57  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_55_sumout ),
	.cout(Xd_0__inst_mult_0_56 ),
	.shareout(Xd_0__inst_mult_0_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_120 (
// Equation(s):
// Xd_0__inst_mult_1_380  = SUM(( GND ) + ( Xd_0__inst_mult_1_378  ) + ( Xd_0__inst_mult_1_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_377 ),
	.sharein(Xd_0__inst_mult_1_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_59 (
// Equation(s):
// Xd_0__inst_mult_1_59_sumout  = SUM(( (din_a[22] & din_b[22]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_60  = CARRY(( (din_a[22] & din_b[22]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_61  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_59_sumout ),
	.cout(Xd_0__inst_mult_1_60 ),
	.shareout(Xd_0__inst_mult_1_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_118 (
// Equation(s):
// Xd_0__inst_mult_9_384  = SUM(( (!din_a[117] & (((din_a[116] & din_b[112])))) # (din_a[117] & (!din_b[111] $ (((!din_a[116]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_486  ) + ( Xd_0__inst_mult_9_485  ))
// Xd_0__inst_mult_9_385  = CARRY(( (!din_a[117] & (((din_a[116] & din_b[112])))) # (din_a[117] & (!din_b[111] $ (((!din_a[116]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_486  ) + ( Xd_0__inst_mult_9_485  ))
// Xd_0__inst_mult_9_386  = SHARE((din_a[117] & (din_b[111] & (din_a[116] & din_b[112]))))

	.dataa(!din_a[117]),
	.datab(!din_b[111]),
	.datac(!din_a[116]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_485 ),
	.sharein(Xd_0__inst_mult_9_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_384 ),
	.cout(Xd_0__inst_mult_9_385 ),
	.shareout(Xd_0__inst_mult_9_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_119 (
// Equation(s):
// Xd_0__inst_mult_9_388  = SUM(( GND ) + ( Xd_0__inst_mult_9_482  ) + ( Xd_0__inst_mult_9_481  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_481 ),
	.sharein(Xd_0__inst_mult_9_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_388 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_118 (
// Equation(s):
// Xd_0__inst_mult_6_384  = SUM(( (!din_a[81] & (((din_a[80] & din_b[76])))) # (din_a[81] & (!din_b[75] $ (((!din_a[80]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_486  ) + ( Xd_0__inst_mult_6_485  ))
// Xd_0__inst_mult_6_385  = CARRY(( (!din_a[81] & (((din_a[80] & din_b[76])))) # (din_a[81] & (!din_b[75] $ (((!din_a[80]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_486  ) + ( Xd_0__inst_mult_6_485  ))
// Xd_0__inst_mult_6_386  = SHARE((din_a[81] & (din_b[75] & (din_a[80] & din_b[76]))))

	.dataa(!din_a[81]),
	.datab(!din_b[75]),
	.datac(!din_a[80]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_485 ),
	.sharein(Xd_0__inst_mult_6_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_384 ),
	.cout(Xd_0__inst_mult_6_385 ),
	.shareout(Xd_0__inst_mult_6_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_119 (
// Equation(s):
// Xd_0__inst_mult_6_388  = SUM(( GND ) + ( Xd_0__inst_mult_6_482  ) + ( Xd_0__inst_mult_6_481  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_481 ),
	.sharein(Xd_0__inst_mult_6_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_388 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_126 (
// Equation(s):
// Xd_0__inst_mult_14_404  = SUM(( (!din_a[175] & (((din_a[174] & din_b[172])))) # (din_a[175] & (!din_b[171] $ (((!din_a[174]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_470  ) + ( Xd_0__inst_mult_14_469  ))
// Xd_0__inst_mult_14_405  = CARRY(( (!din_a[175] & (((din_a[174] & din_b[172])))) # (din_a[175] & (!din_b[171] $ (((!din_a[174]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_470  ) + ( Xd_0__inst_mult_14_469  ))
// Xd_0__inst_mult_14_406  = SHARE((din_a[175] & (din_b[171] & (din_a[174] & din_b[172]))))

	.dataa(!din_a[175]),
	.datab(!din_b[171]),
	.datac(!din_a[174]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_469 ),
	.sharein(Xd_0__inst_mult_14_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_404 ),
	.cout(Xd_0__inst_mult_14_405 ),
	.shareout(Xd_0__inst_mult_14_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_127 (
// Equation(s):
// Xd_0__inst_mult_14_408  = SUM(( (din_a[176] & din_b[170]) ) + ( Xd_0__inst_mult_14_466  ) + ( Xd_0__inst_mult_14_465  ))
// Xd_0__inst_mult_14_409  = CARRY(( (din_a[176] & din_b[170]) ) + ( Xd_0__inst_mult_14_466  ) + ( Xd_0__inst_mult_14_465  ))
// Xd_0__inst_mult_14_410  = SHARE((din_a[178] & din_b[169]))

	.dataa(!din_a[176]),
	.datab(!din_b[170]),
	.datac(!din_a[178]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_465 ),
	.sharein(Xd_0__inst_mult_14_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_408 ),
	.cout(Xd_0__inst_mult_14_409 ),
	.shareout(Xd_0__inst_mult_14_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_122 (
// Equation(s):
// Xd_0__inst_mult_8_388  = SUM(( (!din_a[105] & (((din_a[104] & din_b[100])))) # (din_a[105] & (!din_b[99] $ (((!din_a[104]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_490  ) + ( Xd_0__inst_mult_8_489  ))
// Xd_0__inst_mult_8_389  = CARRY(( (!din_a[105] & (((din_a[104] & din_b[100])))) # (din_a[105] & (!din_b[99] $ (((!din_a[104]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_490  ) + ( Xd_0__inst_mult_8_489  ))
// Xd_0__inst_mult_8_390  = SHARE((din_a[105] & (din_b[99] & (din_a[104] & din_b[100]))))

	.dataa(!din_a[105]),
	.datab(!din_b[99]),
	.datac(!din_a[104]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_489 ),
	.sharein(Xd_0__inst_mult_8_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_388 ),
	.cout(Xd_0__inst_mult_8_389 ),
	.shareout(Xd_0__inst_mult_8_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_123 (
// Equation(s):
// Xd_0__inst_mult_8_392  = SUM(( GND ) + ( Xd_0__inst_mult_8_486  ) + ( Xd_0__inst_mult_8_485  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_485 ),
	.sharein(Xd_0__inst_mult_8_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_392 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_122 (
// Equation(s):
// Xd_0__inst_mult_11_388  = SUM(( (!din_a[141] & (((din_a[140] & din_b[136])))) # (din_a[141] & (!din_b[135] $ (((!din_a[140]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_490  ) + ( Xd_0__inst_mult_11_489  ))
// Xd_0__inst_mult_11_389  = CARRY(( (!din_a[141] & (((din_a[140] & din_b[136])))) # (din_a[141] & (!din_b[135] $ (((!din_a[140]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_490  ) + ( Xd_0__inst_mult_11_489  ))
// Xd_0__inst_mult_11_390  = SHARE((din_a[141] & (din_b[135] & (din_a[140] & din_b[136]))))

	.dataa(!din_a[141]),
	.datab(!din_b[135]),
	.datac(!din_a[140]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_489 ),
	.sharein(Xd_0__inst_mult_11_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_388 ),
	.cout(Xd_0__inst_mult_11_389 ),
	.shareout(Xd_0__inst_mult_11_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_123 (
// Equation(s):
// Xd_0__inst_mult_11_392  = SUM(( GND ) + ( Xd_0__inst_mult_11_486  ) + ( Xd_0__inst_mult_11_485  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_485 ),
	.sharein(Xd_0__inst_mult_11_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_392 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_118 (
// Equation(s):
// Xd_0__inst_mult_10_384  = SUM(( (!din_a[129] & (((din_a[128] & din_b[124])))) # (din_a[129] & (!din_b[123] $ (((!din_a[128]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_486  ) + ( Xd_0__inst_mult_10_485  ))
// Xd_0__inst_mult_10_385  = CARRY(( (!din_a[129] & (((din_a[128] & din_b[124])))) # (din_a[129] & (!din_b[123] $ (((!din_a[128]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_486  ) + ( Xd_0__inst_mult_10_485  ))
// Xd_0__inst_mult_10_386  = SHARE((din_a[129] & (din_b[123] & (din_a[128] & din_b[124]))))

	.dataa(!din_a[129]),
	.datab(!din_b[123]),
	.datac(!din_a[128]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_485 ),
	.sharein(Xd_0__inst_mult_10_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_384 ),
	.cout(Xd_0__inst_mult_10_385 ),
	.shareout(Xd_0__inst_mult_10_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_119 (
// Equation(s):
// Xd_0__inst_mult_10_388  = SUM(( GND ) + ( Xd_0__inst_mult_10_482  ) + ( Xd_0__inst_mult_10_481  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_481 ),
	.sharein(Xd_0__inst_mult_10_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_388 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_128 (
// Equation(s):
// Xd_0__inst_mult_15_412  = SUM(( (din_a[184] & din_b[189]) ) + ( Xd_0__inst_mult_15_538  ) + ( Xd_0__inst_mult_15_537  ))
// Xd_0__inst_mult_15_413  = CARRY(( (din_a[184] & din_b[189]) ) + ( Xd_0__inst_mult_15_538  ) + ( Xd_0__inst_mult_15_537  ))
// Xd_0__inst_mult_15_414  = SHARE((din_a[184] & din_b[190]))

	.dataa(!din_a[184]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_537 ),
	.sharein(Xd_0__inst_mult_15_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_412 ),
	.cout(Xd_0__inst_mult_15_413 ),
	.shareout(Xd_0__inst_mult_15_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_122 (
// Equation(s):
// Xd_0__inst_mult_13_388  = SUM(( (!din_a[165] & (((din_a[164] & din_b[160])))) # (din_a[165] & (!din_b[159] $ (((!din_a[164]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_490  ) + ( Xd_0__inst_mult_13_489  ))
// Xd_0__inst_mult_13_389  = CARRY(( (!din_a[165] & (((din_a[164] & din_b[160])))) # (din_a[165] & (!din_b[159] $ (((!din_a[164]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_490  ) + ( Xd_0__inst_mult_13_489  ))
// Xd_0__inst_mult_13_390  = SHARE((din_a[165] & (din_b[159] & (din_a[164] & din_b[160]))))

	.dataa(!din_a[165]),
	.datab(!din_b[159]),
	.datac(!din_a[164]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_489 ),
	.sharein(Xd_0__inst_mult_13_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_388 ),
	.cout(Xd_0__inst_mult_13_389 ),
	.shareout(Xd_0__inst_mult_13_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_123 (
// Equation(s):
// Xd_0__inst_mult_13_392  = SUM(( GND ) + ( Xd_0__inst_mult_13_486  ) + ( Xd_0__inst_mult_13_485  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_485 ),
	.sharein(Xd_0__inst_mult_13_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_392 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_129 (
// Equation(s):
// Xd_0__inst_mult_15_416  = SUM(( (!din_a[189] & (((din_a[188] & din_b[184])))) # (din_a[189] & (!din_b[183] $ (((!din_a[188]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_518  ) + ( Xd_0__inst_mult_15_517  ))
// Xd_0__inst_mult_15_417  = CARRY(( (!din_a[189] & (((din_a[188] & din_b[184])))) # (din_a[189] & (!din_b[183] $ (((!din_a[188]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_518  ) + ( Xd_0__inst_mult_15_517  ))
// Xd_0__inst_mult_15_418  = SHARE((din_a[189] & (din_b[183] & (din_a[188] & din_b[184]))))

	.dataa(!din_a[189]),
	.datab(!din_b[183]),
	.datac(!din_a[188]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_517 ),
	.sharein(Xd_0__inst_mult_15_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_416 ),
	.cout(Xd_0__inst_mult_15_417 ),
	.shareout(Xd_0__inst_mult_15_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_130 (
// Equation(s):
// Xd_0__inst_mult_15_420  = SUM(( GND ) + ( Xd_0__inst_mult_15_514  ) + ( Xd_0__inst_mult_15_513  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_513 ),
	.sharein(Xd_0__inst_mult_15_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_420 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_124 (
// Equation(s):
// Xd_0__inst_mult_12_408  = SUM(( (!din_a[153] & (((din_a[152] & din_b[148])))) # (din_a[153] & (!din_b[147] $ (((!din_a[152]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_514  ) + ( Xd_0__inst_mult_12_513  ))
// Xd_0__inst_mult_12_409  = CARRY(( (!din_a[153] & (((din_a[152] & din_b[148])))) # (din_a[153] & (!din_b[147] $ (((!din_a[152]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_514  ) + ( Xd_0__inst_mult_12_513  ))
// Xd_0__inst_mult_12_410  = SHARE((din_a[153] & (din_b[147] & (din_a[152] & din_b[148]))))

	.dataa(!din_a[153]),
	.datab(!din_b[147]),
	.datac(!din_a[152]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_513 ),
	.sharein(Xd_0__inst_mult_12_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_408 ),
	.cout(Xd_0__inst_mult_12_409 ),
	.shareout(Xd_0__inst_mult_12_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_125 (
// Equation(s):
// Xd_0__inst_mult_12_412  = SUM(( GND ) + ( Xd_0__inst_mult_12_510  ) + ( Xd_0__inst_mult_12_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_509 ),
	.sharein(Xd_0__inst_mult_12_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_412 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_126 (
// Equation(s):
// Xd_0__inst_mult_12_416  = SUM(( (din_a[148] & din_b[153]) ) + ( Xd_0__inst_mult_12_534  ) + ( Xd_0__inst_mult_12_533  ))
// Xd_0__inst_mult_12_417  = CARRY(( (din_a[148] & din_b[153]) ) + ( Xd_0__inst_mult_12_534  ) + ( Xd_0__inst_mult_12_533  ))
// Xd_0__inst_mult_12_418  = SHARE((din_a[148] & din_b[154]))

	.dataa(!din_a[148]),
	.datab(!din_b[153]),
	.datac(!din_b[154]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_533 ),
	.sharein(Xd_0__inst_mult_12_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_416 ),
	.cout(Xd_0__inst_mult_12_417 ),
	.shareout(Xd_0__inst_mult_12_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_128 (
// Equation(s):
// Xd_0__inst_mult_4_412  = SUM(( (din_a[50] & din_b[57]) ) + ( Xd_0__inst_mult_4_498  ) + ( Xd_0__inst_mult_4_497  ))
// Xd_0__inst_mult_4_413  = CARRY(( (din_a[50] & din_b[57]) ) + ( Xd_0__inst_mult_4_498  ) + ( Xd_0__inst_mult_4_497  ))
// Xd_0__inst_mult_4_414  = SHARE((din_a[50] & din_b[58]))

	.dataa(!din_a[50]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_497 ),
	.sharein(Xd_0__inst_mult_4_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_412 ),
	.cout(Xd_0__inst_mult_4_413 ),
	.shareout(Xd_0__inst_mult_4_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_127 (
// Equation(s):
// Xd_0__inst_mult_12_420  = SUM(( (!din_a[146] & (((din_a[147] & din_b[144])))) # (din_a[146] & (!din_b[145] $ (((!din_a[147]) # (!din_b[144]))))) ) + ( Xd_0__inst_mult_12_282  ) + ( Xd_0__inst_mult_12_281  ))
// Xd_0__inst_mult_12_421  = CARRY(( (!din_a[146] & (((din_a[147] & din_b[144])))) # (din_a[146] & (!din_b[145] $ (((!din_a[147]) # (!din_b[144]))))) ) + ( Xd_0__inst_mult_12_282  ) + ( Xd_0__inst_mult_12_281  ))
// Xd_0__inst_mult_12_422  = SHARE((din_a[146] & (din_b[145] & (din_a[147] & din_b[144]))))

	.dataa(!din_a[146]),
	.datab(!din_b[145]),
	.datac(!din_a[147]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_281 ),
	.sharein(Xd_0__inst_mult_12_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_420 ),
	.cout(Xd_0__inst_mult_12_421 ),
	.shareout(Xd_0__inst_mult_12_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_128 (
// Equation(s):
// Xd_0__inst_mult_12_425  = CARRY(( GND ) + ( Xd_0__inst_mult_13_65  ) + ( Xd_0__inst_mult_13_64  ))
// Xd_0__inst_mult_12_426  = SHARE(Xd_0__inst_mult_12_420 )

	.dataa(!Xd_0__inst_mult_12_420 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_64 ),
	.sharein(Xd_0__inst_mult_13_65 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_425 ),
	.shareout(Xd_0__inst_mult_12_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_124 (
// Equation(s):
// Xd_0__inst_mult_13_396  = SUM(( (!din_a[158] & (((din_a[159] & din_b[156])))) # (din_a[158] & (!din_b[157] $ (((!din_a[159]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_13_266  ) + ( Xd_0__inst_mult_13_265  ))
// Xd_0__inst_mult_13_397  = CARRY(( (!din_a[158] & (((din_a[159] & din_b[156])))) # (din_a[158] & (!din_b[157] $ (((!din_a[159]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_13_266  ) + ( Xd_0__inst_mult_13_265  ))
// Xd_0__inst_mult_13_398  = SHARE((din_a[158] & (din_b[157] & (din_a[159] & din_b[156]))))

	.dataa(!din_a[158]),
	.datab(!din_b[157]),
	.datac(!din_a[159]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_265 ),
	.sharein(Xd_0__inst_mult_13_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_396 ),
	.cout(Xd_0__inst_mult_13_397 ),
	.shareout(Xd_0__inst_mult_13_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_125 (
// Equation(s):
// Xd_0__inst_mult_13_401  = CARRY(( GND ) + ( Xd_0__inst_mult_4_61  ) + ( Xd_0__inst_mult_4_60  ))
// Xd_0__inst_mult_13_402  = SHARE(Xd_0__inst_mult_13_396 )

	.dataa(!Xd_0__inst_mult_13_396 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_60 ),
	.sharein(Xd_0__inst_mult_4_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_401 ),
	.shareout(Xd_0__inst_mult_13_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_128 (
// Equation(s):
// Xd_0__inst_mult_14_412  = SUM(( (!din_a[170] & (((din_a[171] & din_b[168])))) # (din_a[170] & (!din_b[169] $ (((!din_a[171]) # (!din_b[168]))))) ) + ( Xd_0__inst_mult_14_286  ) + ( Xd_0__inst_mult_14_285  ))
// Xd_0__inst_mult_14_413  = CARRY(( (!din_a[170] & (((din_a[171] & din_b[168])))) # (din_a[170] & (!din_b[169] $ (((!din_a[171]) # (!din_b[168]))))) ) + ( Xd_0__inst_mult_14_286  ) + ( Xd_0__inst_mult_14_285  ))
// Xd_0__inst_mult_14_414  = SHARE((din_a[170] & (din_b[169] & (din_a[171] & din_b[168]))))

	.dataa(!din_a[170]),
	.datab(!din_b[169]),
	.datac(!din_a[171]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_285 ),
	.sharein(Xd_0__inst_mult_14_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_412 ),
	.cout(Xd_0__inst_mult_14_413 ),
	.shareout(Xd_0__inst_mult_14_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_129 (
// Equation(s):
// Xd_0__inst_mult_14_417  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_418  = SHARE(Xd_0__inst_mult_14_412 )

	.dataa(!Xd_0__inst_mult_14_412 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_417 ),
	.shareout(Xd_0__inst_mult_14_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_131 (
// Equation(s):
// Xd_0__inst_mult_15_424  = SUM(( (!din_a[182] & (((din_a[183] & din_b[180])))) # (din_a[182] & (!din_b[181] $ (((!din_a[183]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_15_286  ) + ( Xd_0__inst_mult_15_285  ))
// Xd_0__inst_mult_15_425  = CARRY(( (!din_a[182] & (((din_a[183] & din_b[180])))) # (din_a[182] & (!din_b[181] $ (((!din_a[183]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_15_286  ) + ( Xd_0__inst_mult_15_285  ))
// Xd_0__inst_mult_15_426  = SHARE((din_a[182] & (din_b[181] & (din_a[183] & din_b[180]))))

	.dataa(!din_a[182]),
	.datab(!din_b[181]),
	.datac(!din_a[183]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_285 ),
	.sharein(Xd_0__inst_mult_15_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_424 ),
	.cout(Xd_0__inst_mult_15_425 ),
	.shareout(Xd_0__inst_mult_15_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_132 (
// Equation(s):
// Xd_0__inst_mult_15_429  = CARRY(( GND ) + ( Xd_0__inst_mult_5_61  ) + ( Xd_0__inst_mult_5_60  ))
// Xd_0__inst_mult_15_430  = SHARE(Xd_0__inst_mult_15_424 )

	.dataa(!Xd_0__inst_mult_15_424 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_60 ),
	.sharein(Xd_0__inst_mult_5_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_429 ),
	.shareout(Xd_0__inst_mult_15_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_120 (
// Equation(s):
// Xd_0__inst_mult_10_392  = SUM(( (!din_a[122] & (((din_a[123] & din_b[120])))) # (din_a[122] & (!din_b[121] $ (((!din_a[123]) # (!din_b[120]))))) ) + ( Xd_0__inst_mult_10_262  ) + ( Xd_0__inst_mult_10_261  ))
// Xd_0__inst_mult_10_393  = CARRY(( (!din_a[122] & (((din_a[123] & din_b[120])))) # (din_a[122] & (!din_b[121] $ (((!din_a[123]) # (!din_b[120]))))) ) + ( Xd_0__inst_mult_10_262  ) + ( Xd_0__inst_mult_10_261  ))
// Xd_0__inst_mult_10_394  = SHARE((din_a[122] & (din_b[121] & (din_a[123] & din_b[120]))))

	.dataa(!din_a[122]),
	.datab(!din_b[121]),
	.datac(!din_a[123]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_261 ),
	.sharein(Xd_0__inst_mult_10_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_392 ),
	.cout(Xd_0__inst_mult_10_393 ),
	.shareout(Xd_0__inst_mult_10_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_121 (
// Equation(s):
// Xd_0__inst_mult_10_397  = CARRY(( GND ) + ( Xd_0__inst_mult_7_57  ) + ( Xd_0__inst_mult_7_56  ))
// Xd_0__inst_mult_10_398  = SHARE(Xd_0__inst_mult_10_392 )

	.dataa(!Xd_0__inst_mult_10_392 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_56 ),
	.sharein(Xd_0__inst_mult_7_57 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_397 ),
	.shareout(Xd_0__inst_mult_10_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_124 (
// Equation(s):
// Xd_0__inst_mult_11_396  = SUM(( (!din_a[134] & (((din_a[135] & din_b[132])))) # (din_a[134] & (!din_b[133] $ (((!din_a[135]) # (!din_b[132]))))) ) + ( Xd_0__inst_mult_11_266  ) + ( Xd_0__inst_mult_11_265  ))
// Xd_0__inst_mult_11_397  = CARRY(( (!din_a[134] & (((din_a[135] & din_b[132])))) # (din_a[134] & (!din_b[133] $ (((!din_a[135]) # (!din_b[132]))))) ) + ( Xd_0__inst_mult_11_266  ) + ( Xd_0__inst_mult_11_265  ))
// Xd_0__inst_mult_11_398  = SHARE((din_a[134] & (din_b[133] & (din_a[135] & din_b[132]))))

	.dataa(!din_a[134]),
	.datab(!din_b[133]),
	.datac(!din_a[135]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_265 ),
	.sharein(Xd_0__inst_mult_11_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_396 ),
	.cout(Xd_0__inst_mult_11_397 ),
	.shareout(Xd_0__inst_mult_11_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_125 (
// Equation(s):
// Xd_0__inst_mult_11_401  = CARRY(( GND ) + ( Xd_0__inst_mult_6_61  ) + ( Xd_0__inst_mult_6_60  ))
// Xd_0__inst_mult_11_402  = SHARE(Xd_0__inst_mult_11_396 )

	.dataa(!Xd_0__inst_mult_11_396 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_60 ),
	.sharein(Xd_0__inst_mult_6_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_401 ),
	.shareout(Xd_0__inst_mult_11_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_124 (
// Equation(s):
// Xd_0__inst_mult_8_396  = SUM(( (!din_a[98] & (((din_a[99] & din_b[96])))) # (din_a[98] & (!din_b[97] $ (((!din_a[99]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_8_266  ) + ( Xd_0__inst_mult_8_265  ))
// Xd_0__inst_mult_8_397  = CARRY(( (!din_a[98] & (((din_a[99] & din_b[96])))) # (din_a[98] & (!din_b[97] $ (((!din_a[99]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_8_266  ) + ( Xd_0__inst_mult_8_265  ))
// Xd_0__inst_mult_8_398  = SHARE((din_a[98] & (din_b[97] & (din_a[99] & din_b[96]))))

	.dataa(!din_a[98]),
	.datab(!din_b[97]),
	.datac(!din_a[99]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_265 ),
	.sharein(Xd_0__inst_mult_8_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_396 ),
	.cout(Xd_0__inst_mult_8_397 ),
	.shareout(Xd_0__inst_mult_8_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_125 (
// Equation(s):
// Xd_0__inst_mult_8_401  = CARRY(( GND ) + ( Xd_0__inst_mult_9_61  ) + ( Xd_0__inst_mult_9_60  ))
// Xd_0__inst_mult_8_402  = SHARE(Xd_0__inst_mult_8_396 )

	.dataa(!Xd_0__inst_mult_8_396 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_60 ),
	.sharein(Xd_0__inst_mult_9_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_401 ),
	.shareout(Xd_0__inst_mult_8_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_120 (
// Equation(s):
// Xd_0__inst_mult_9_392  = SUM(( (!din_a[110] & (((din_a[111] & din_b[108])))) # (din_a[110] & (!din_b[109] $ (((!din_a[111]) # (!din_b[108]))))) ) + ( Xd_0__inst_mult_9_262  ) + ( Xd_0__inst_mult_9_261  ))
// Xd_0__inst_mult_9_393  = CARRY(( (!din_a[110] & (((din_a[111] & din_b[108])))) # (din_a[110] & (!din_b[109] $ (((!din_a[111]) # (!din_b[108]))))) ) + ( Xd_0__inst_mult_9_262  ) + ( Xd_0__inst_mult_9_261  ))
// Xd_0__inst_mult_9_394  = SHARE((din_a[110] & (din_b[109] & (din_a[111] & din_b[108]))))

	.dataa(!din_a[110]),
	.datab(!din_b[109]),
	.datac(!din_a[111]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_261 ),
	.sharein(Xd_0__inst_mult_9_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_392 ),
	.cout(Xd_0__inst_mult_9_393 ),
	.shareout(Xd_0__inst_mult_9_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_121 (
// Equation(s):
// Xd_0__inst_mult_9_397  = CARRY(( GND ) + ( Xd_0__inst_mult_8_65  ) + ( Xd_0__inst_mult_8_64  ))
// Xd_0__inst_mult_9_398  = SHARE(Xd_0__inst_mult_9_392 )

	.dataa(!Xd_0__inst_mult_9_392 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_64 ),
	.sharein(Xd_0__inst_mult_8_65 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_397 ),
	.shareout(Xd_0__inst_mult_9_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_120 (
// Equation(s):
// Xd_0__inst_mult_6_392  = SUM(( (!din_a[74] & (((din_a[75] & din_b[72])))) # (din_a[74] & (!din_b[73] $ (((!din_a[75]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_262  ) + ( Xd_0__inst_mult_6_261  ))
// Xd_0__inst_mult_6_393  = CARRY(( (!din_a[74] & (((din_a[75] & din_b[72])))) # (din_a[74] & (!din_b[73] $ (((!din_a[75]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_262  ) + ( Xd_0__inst_mult_6_261  ))
// Xd_0__inst_mult_6_394  = SHARE((din_a[74] & (din_b[73] & (din_a[75] & din_b[72]))))

	.dataa(!din_a[74]),
	.datab(!din_b[73]),
	.datac(!din_a[75]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_261 ),
	.sharein(Xd_0__inst_mult_6_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_392 ),
	.cout(Xd_0__inst_mult_6_393 ),
	.shareout(Xd_0__inst_mult_6_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_121 (
// Equation(s):
// Xd_0__inst_mult_6_397  = CARRY(( GND ) + ( Xd_0__inst_mult_11_65  ) + ( Xd_0__inst_mult_11_64  ))
// Xd_0__inst_mult_6_398  = SHARE(Xd_0__inst_mult_6_392 )

	.dataa(!Xd_0__inst_mult_6_392 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_64 ),
	.sharein(Xd_0__inst_mult_11_65 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_397 ),
	.shareout(Xd_0__inst_mult_6_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_116 (
// Equation(s):
// Xd_0__inst_mult_7_376  = SUM(( (!din_a[86] & (((din_a[87] & din_b[84])))) # (din_a[86] & (!din_b[85] $ (((!din_a[87]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_246  ) + ( Xd_0__inst_mult_7_245  ))
// Xd_0__inst_mult_7_377  = CARRY(( (!din_a[86] & (((din_a[87] & din_b[84])))) # (din_a[86] & (!din_b[85] $ (((!din_a[87]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_246  ) + ( Xd_0__inst_mult_7_245  ))
// Xd_0__inst_mult_7_378  = SHARE((din_a[86] & (din_b[85] & (din_a[87] & din_b[84]))))

	.dataa(!din_a[86]),
	.datab(!din_b[85]),
	.datac(!din_a[87]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_245 ),
	.sharein(Xd_0__inst_mult_7_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_376 ),
	.cout(Xd_0__inst_mult_7_377 ),
	.shareout(Xd_0__inst_mult_7_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_117 (
// Equation(s):
// Xd_0__inst_mult_7_380  = SUM(( (din_a[70] & din_b[60]) ) + ( Xd_0__inst_mult_2_69  ) + ( Xd_0__inst_mult_2_68  ))
// Xd_0__inst_mult_7_381  = CARRY(( (din_a[70] & din_b[60]) ) + ( Xd_0__inst_mult_2_69  ) + ( Xd_0__inst_mult_2_68  ))
// Xd_0__inst_mult_7_382  = SHARE(Xd_0__inst_mult_7_376 )

	.dataa(!din_a[70]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_7_376 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_68 ),
	.sharein(Xd_0__inst_mult_2_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_380 ),
	.cout(Xd_0__inst_mult_7_381 ),
	.shareout(Xd_0__inst_mult_7_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_129 (
// Equation(s):
// Xd_0__inst_mult_4_416  = SUM(( (!din_a[50] & (((din_a[51] & din_b[48])))) # (din_a[50] & (!din_b[49] $ (((!din_a[51]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_278  ) + ( Xd_0__inst_mult_4_277  ))
// Xd_0__inst_mult_4_417  = CARRY(( (!din_a[50] & (((din_a[51] & din_b[48])))) # (din_a[50] & (!din_b[49] $ (((!din_a[51]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_278  ) + ( Xd_0__inst_mult_4_277  ))
// Xd_0__inst_mult_4_418  = SHARE((din_a[50] & (din_b[49] & (din_a[51] & din_b[48]))))

	.dataa(!din_a[50]),
	.datab(!din_b[49]),
	.datac(!din_a[51]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_277 ),
	.sharein(Xd_0__inst_mult_4_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_416 ),
	.cout(Xd_0__inst_mult_4_417 ),
	.shareout(Xd_0__inst_mult_4_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_130 (
// Equation(s):
// Xd_0__inst_mult_4_420  = SUM(( (din_a[80] & din_b[72]) ) + ( Xd_0__inst_mult_7_61  ) + ( Xd_0__inst_mult_7_60  ))
// Xd_0__inst_mult_4_421  = CARRY(( (din_a[80] & din_b[72]) ) + ( Xd_0__inst_mult_7_61  ) + ( Xd_0__inst_mult_7_60  ))
// Xd_0__inst_mult_4_422  = SHARE(Xd_0__inst_mult_4_416 )

	.dataa(!din_a[80]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_4_416 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_60 ),
	.sharein(Xd_0__inst_mult_7_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_420 ),
	.cout(Xd_0__inst_mult_4_421 ),
	.shareout(Xd_0__inst_mult_4_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_116 (
// Equation(s):
// Xd_0__inst_mult_5_376  = SUM(( (!din_a[62] & (((din_a[63] & din_b[60])))) # (din_a[62] & (!din_b[61] $ (((!din_a[63]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_246  ) + ( Xd_0__inst_mult_5_245  ))
// Xd_0__inst_mult_5_377  = CARRY(( (!din_a[62] & (((din_a[63] & din_b[60])))) # (din_a[62] & (!din_b[61] $ (((!din_a[63]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_246  ) + ( Xd_0__inst_mult_5_245  ))
// Xd_0__inst_mult_5_378  = SHARE((din_a[62] & (din_b[61] & (din_a[63] & din_b[60]))))

	.dataa(!din_a[62]),
	.datab(!din_b[61]),
	.datac(!din_a[63]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_245 ),
	.sharein(Xd_0__inst_mult_5_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_376 ),
	.cout(Xd_0__inst_mult_5_377 ),
	.shareout(Xd_0__inst_mult_5_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_117 (
// Equation(s):
// Xd_0__inst_mult_5_380  = SUM(( (din_a[44] & din_b[36]) ) + ( Xd_0__inst_mult_0_65  ) + ( Xd_0__inst_mult_0_64  ))
// Xd_0__inst_mult_5_381  = CARRY(( (din_a[44] & din_b[36]) ) + ( Xd_0__inst_mult_0_65  ) + ( Xd_0__inst_mult_0_64  ))
// Xd_0__inst_mult_5_382  = SHARE(Xd_0__inst_mult_5_376 )

	.dataa(!din_a[44]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_5_376 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_64 ),
	.sharein(Xd_0__inst_mult_0_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_380 ),
	.cout(Xd_0__inst_mult_5_381 ),
	.shareout(Xd_0__inst_mult_5_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_120 (
// Equation(s):
// Xd_0__inst_mult_2_380  = SUM(( (!din_a[26] & (((din_a[27] & din_b[24])))) # (din_a[26] & (!din_b[25] $ (((!din_a[27]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_250  ) + ( Xd_0__inst_mult_2_249  ))
// Xd_0__inst_mult_2_381  = CARRY(( (!din_a[26] & (((din_a[27] & din_b[24])))) # (din_a[26] & (!din_b[25] $ (((!din_a[27]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_250  ) + ( Xd_0__inst_mult_2_249  ))
// Xd_0__inst_mult_2_382  = SHARE((din_a[26] & (din_b[25] & (din_a[27] & din_b[24]))))

	.dataa(!din_a[26]),
	.datab(!din_b[25]),
	.datac(!din_a[27]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_249 ),
	.sharein(Xd_0__inst_mult_2_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_380 ),
	.cout(Xd_0__inst_mult_2_381 ),
	.shareout(Xd_0__inst_mult_2_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_121 (
// Equation(s):
// Xd_0__inst_mult_2_384  = SUM(( (din_a[153] & din_b[144]) ) + ( Xd_0__inst_mult_13_69  ) + ( Xd_0__inst_mult_13_68  ))
// Xd_0__inst_mult_2_385  = CARRY(( (din_a[153] & din_b[144]) ) + ( Xd_0__inst_mult_13_69  ) + ( Xd_0__inst_mult_13_68  ))
// Xd_0__inst_mult_2_386  = SHARE(Xd_0__inst_mult_2_380 )

	.dataa(!din_a[153]),
	.datab(!din_b[144]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_2_380 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_68 ),
	.sharein(Xd_0__inst_mult_13_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_384 ),
	.cout(Xd_0__inst_mult_2_385 ),
	.shareout(Xd_0__inst_mult_2_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_116 (
// Equation(s):
// Xd_0__inst_mult_3_376  = SUM(( (!din_a[38] & (((din_a[39] & din_b[36])))) # (din_a[38] & (!din_b[37] $ (((!din_a[39]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_246  ) + ( Xd_0__inst_mult_3_245  ))
// Xd_0__inst_mult_3_377  = CARRY(( (!din_a[38] & (((din_a[39] & din_b[36])))) # (din_a[38] & (!din_b[37] $ (((!din_a[39]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_246  ) + ( Xd_0__inst_mult_3_245  ))
// Xd_0__inst_mult_3_378  = SHARE((din_a[38] & (din_b[37] & (din_a[39] & din_b[36]))))

	.dataa(!din_a[38]),
	.datab(!din_b[37]),
	.datac(!din_a[39]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_245 ),
	.sharein(Xd_0__inst_mult_3_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_376 ),
	.cout(Xd_0__inst_mult_3_377 ),
	.shareout(Xd_0__inst_mult_3_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_117 (
// Equation(s):
// Xd_0__inst_mult_3_380  = SUM(( (din_a[117] & din_b[108]) ) + ( Xd_0__inst_mult_6_65  ) + ( Xd_0__inst_mult_6_64  ))
// Xd_0__inst_mult_3_381  = CARRY(( (din_a[117] & din_b[108]) ) + ( Xd_0__inst_mult_6_65  ) + ( Xd_0__inst_mult_6_64  ))
// Xd_0__inst_mult_3_382  = SHARE(Xd_0__inst_mult_3_376 )

	.dataa(!din_a[117]),
	.datab(!din_b[108]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_3_376 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_64 ),
	.sharein(Xd_0__inst_mult_6_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_380 ),
	.cout(Xd_0__inst_mult_3_381 ),
	.shareout(Xd_0__inst_mult_3_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_121 (
// Equation(s):
// Xd_0__inst_mult_0_384  = SUM(( (!din_a[2] & (((din_a[3] & din_b[0])))) # (din_a[2] & (!din_b[1] $ (((!din_a[3]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_250  ) + ( Xd_0__inst_mult_0_249  ))
// Xd_0__inst_mult_0_385  = CARRY(( (!din_a[2] & (((din_a[3] & din_b[0])))) # (din_a[2] & (!din_b[1] $ (((!din_a[3]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_250  ) + ( Xd_0__inst_mult_0_249  ))
// Xd_0__inst_mult_0_386  = SHARE((din_a[2] & (din_b[1] & (din_a[3] & din_b[0]))))

	.dataa(!din_a[2]),
	.datab(!din_b[1]),
	.datac(!din_a[3]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_249 ),
	.sharein(Xd_0__inst_mult_0_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_384 ),
	.cout(Xd_0__inst_mult_0_385 ),
	.shareout(Xd_0__inst_mult_0_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_121 (
// Equation(s):
// Xd_0__inst_mult_1_384  = SUM(( (!din_a[14] & (((din_a[15] & din_b[12])))) # (din_a[14] & (!din_b[13] $ (((!din_a[15]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_250  ) + ( Xd_0__inst_mult_1_249  ))
// Xd_0__inst_mult_1_385  = CARRY(( (!din_a[14] & (((din_a[15] & din_b[12])))) # (din_a[14] & (!din_b[13] $ (((!din_a[15]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_250  ) + ( Xd_0__inst_mult_1_249  ))
// Xd_0__inst_mult_1_386  = SHARE((din_a[14] & (din_b[13] & (din_a[15] & din_b[12]))))

	.dataa(!din_a[14]),
	.datab(!din_b[13]),
	.datac(!din_a[15]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_249 ),
	.sharein(Xd_0__inst_mult_1_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_384 ),
	.cout(Xd_0__inst_mult_1_385 ),
	.shareout(Xd_0__inst_mult_1_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_129 (
// Equation(s):
// Xd_0__inst_mult_12_429  = CARRY(( (din_a[147] & din_b[145]) ) + ( Xd_0__inst_mult_12_570  ) + ( Xd_0__inst_mult_12_569  ))
// Xd_0__inst_mult_12_430  = SHARE((din_a[146] & din_b[146]))

	.dataa(!din_a[147]),
	.datab(!din_b[145]),
	.datac(!din_a[146]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_569 ),
	.sharein(Xd_0__inst_mult_12_570 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_429 ),
	.shareout(Xd_0__inst_mult_12_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_126 (
// Equation(s):
// Xd_0__inst_mult_13_405  = CARRY(( (din_a[159] & din_b[157]) ) + ( Xd_0__inst_mult_13_578  ) + ( Xd_0__inst_mult_13_577  ))
// Xd_0__inst_mult_13_406  = SHARE((din_a[158] & din_b[158]))

	.dataa(!din_a[159]),
	.datab(!din_b[157]),
	.datac(!din_a[158]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_577 ),
	.sharein(Xd_0__inst_mult_13_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_405 ),
	.shareout(Xd_0__inst_mult_13_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_130 (
// Equation(s):
// Xd_0__inst_mult_14_421  = CARRY(( (din_a[171] & din_b[169]) ) + ( Xd_0__inst_mult_14_554  ) + ( Xd_0__inst_mult_14_553  ))
// Xd_0__inst_mult_14_422  = SHARE((din_a[170] & din_b[170]))

	.dataa(!din_a[171]),
	.datab(!din_b[169]),
	.datac(!din_a[170]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_553 ),
	.sharein(Xd_0__inst_mult_14_554 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_421 ),
	.shareout(Xd_0__inst_mult_14_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_133 (
// Equation(s):
// Xd_0__inst_mult_15_433  = CARRY(( (din_a[183] & din_b[181]) ) + ( Xd_0__inst_mult_15_562  ) + ( Xd_0__inst_mult_15_561  ))
// Xd_0__inst_mult_15_434  = SHARE((din_a[182] & din_b[182]))

	.dataa(!din_a[183]),
	.datab(!din_b[181]),
	.datac(!din_a[182]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_561 ),
	.sharein(Xd_0__inst_mult_15_562 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_433 ),
	.shareout(Xd_0__inst_mult_15_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_122 (
// Equation(s):
// Xd_0__inst_mult_10_401  = CARRY(( (din_a[123] & din_b[121]) ) + ( Xd_0__inst_mult_10_574  ) + ( Xd_0__inst_mult_10_573  ))
// Xd_0__inst_mult_10_402  = SHARE((din_a[122] & din_b[122]))

	.dataa(!din_a[123]),
	.datab(!din_b[121]),
	.datac(!din_a[122]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_573 ),
	.sharein(Xd_0__inst_mult_10_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_401 ),
	.shareout(Xd_0__inst_mult_10_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_126 (
// Equation(s):
// Xd_0__inst_mult_11_405  = CARRY(( (din_a[135] & din_b[133]) ) + ( Xd_0__inst_mult_11_578  ) + ( Xd_0__inst_mult_11_577  ))
// Xd_0__inst_mult_11_406  = SHARE((din_a[134] & din_b[134]))

	.dataa(!din_a[135]),
	.datab(!din_b[133]),
	.datac(!din_a[134]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_577 ),
	.sharein(Xd_0__inst_mult_11_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_405 ),
	.shareout(Xd_0__inst_mult_11_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_126 (
// Equation(s):
// Xd_0__inst_mult_8_405  = CARRY(( (din_a[99] & din_b[97]) ) + ( Xd_0__inst_mult_8_578  ) + ( Xd_0__inst_mult_8_577  ))
// Xd_0__inst_mult_8_406  = SHARE((din_a[98] & din_b[98]))

	.dataa(!din_a[99]),
	.datab(!din_b[97]),
	.datac(!din_a[98]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_577 ),
	.sharein(Xd_0__inst_mult_8_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_405 ),
	.shareout(Xd_0__inst_mult_8_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_122 (
// Equation(s):
// Xd_0__inst_mult_9_401  = CARRY(( (din_a[111] & din_b[109]) ) + ( Xd_0__inst_mult_9_574  ) + ( Xd_0__inst_mult_9_573  ))
// Xd_0__inst_mult_9_402  = SHARE((din_a[110] & din_b[110]))

	.dataa(!din_a[111]),
	.datab(!din_b[109]),
	.datac(!din_a[110]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_573 ),
	.sharein(Xd_0__inst_mult_9_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_401 ),
	.shareout(Xd_0__inst_mult_9_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_122 (
// Equation(s):
// Xd_0__inst_mult_6_401  = CARRY(( (din_a[75] & din_b[73]) ) + ( Xd_0__inst_mult_6_574  ) + ( Xd_0__inst_mult_6_573  ))
// Xd_0__inst_mult_6_402  = SHARE((din_a[74] & din_b[74]))

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_573 ),
	.sharein(Xd_0__inst_mult_6_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_401 ),
	.shareout(Xd_0__inst_mult_6_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_118 (
// Equation(s):
// Xd_0__inst_mult_7_385  = CARRY(( (din_a[87] & din_b[85]) ) + ( Xd_0__inst_mult_7_574  ) + ( Xd_0__inst_mult_7_573  ))
// Xd_0__inst_mult_7_386  = SHARE((din_a[86] & din_b[86]))

	.dataa(!din_a[87]),
	.datab(!din_b[85]),
	.datac(!din_a[86]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_573 ),
	.sharein(Xd_0__inst_mult_7_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_385 ),
	.shareout(Xd_0__inst_mult_7_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_131 (
// Equation(s):
// Xd_0__inst_mult_4_425  = CARRY(( (din_a[51] & din_b[49]) ) + ( Xd_0__inst_mult_4_574  ) + ( Xd_0__inst_mult_4_573  ))
// Xd_0__inst_mult_4_426  = SHARE((din_a[50] & din_b[50]))

	.dataa(!din_a[51]),
	.datab(!din_b[49]),
	.datac(!din_a[50]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_573 ),
	.sharein(Xd_0__inst_mult_4_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_425 ),
	.shareout(Xd_0__inst_mult_4_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_118 (
// Equation(s):
// Xd_0__inst_mult_5_385  = CARRY(( (din_a[63] & din_b[61]) ) + ( Xd_0__inst_mult_5_574  ) + ( Xd_0__inst_mult_5_573  ))
// Xd_0__inst_mult_5_386  = SHARE((din_a[62] & din_b[62]))

	.dataa(!din_a[63]),
	.datab(!din_b[61]),
	.datac(!din_a[62]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_573 ),
	.sharein(Xd_0__inst_mult_5_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_385 ),
	.shareout(Xd_0__inst_mult_5_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_122 (
// Equation(s):
// Xd_0__inst_mult_2_389  = CARRY(( (din_a[27] & din_b[25]) ) + ( Xd_0__inst_mult_2_578  ) + ( Xd_0__inst_mult_2_577  ))
// Xd_0__inst_mult_2_390  = SHARE((din_a[26] & din_b[26]))

	.dataa(!din_a[27]),
	.datab(!din_b[25]),
	.datac(!din_a[26]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_577 ),
	.sharein(Xd_0__inst_mult_2_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_389 ),
	.shareout(Xd_0__inst_mult_2_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_118 (
// Equation(s):
// Xd_0__inst_mult_3_385  = CARRY(( (din_a[39] & din_b[37]) ) + ( Xd_0__inst_mult_3_574  ) + ( Xd_0__inst_mult_3_573  ))
// Xd_0__inst_mult_3_386  = SHARE((din_a[38] & din_b[38]))

	.dataa(!din_a[39]),
	.datab(!din_b[37]),
	.datac(!din_a[38]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_573 ),
	.sharein(Xd_0__inst_mult_3_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_385 ),
	.shareout(Xd_0__inst_mult_3_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_122 (
// Equation(s):
// Xd_0__inst_mult_0_389  = CARRY(( (din_a[3] & din_b[1]) ) + ( Xd_0__inst_mult_0_578  ) + ( Xd_0__inst_mult_0_577  ))
// Xd_0__inst_mult_0_390  = SHARE((din_a[2] & din_b[2]))

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_577 ),
	.sharein(Xd_0__inst_mult_0_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_389 ),
	.shareout(Xd_0__inst_mult_0_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_122 (
// Equation(s):
// Xd_0__inst_mult_1_389  = CARRY(( (din_a[15] & din_b[13]) ) + ( Xd_0__inst_mult_1_542  ) + ( Xd_0__inst_mult_1_541  ))
// Xd_0__inst_mult_1_390  = SHARE((din_a[14] & din_b[14]))

	.dataa(!din_a[15]),
	.datab(!din_b[13]),
	.datac(!din_a[14]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_541 ),
	.sharein(Xd_0__inst_mult_1_542 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_389 ),
	.shareout(Xd_0__inst_mult_1_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_130 (
// Equation(s):
// Xd_0__inst_mult_12_432  = SUM(( (din_a[149] & din_b[144]) ) + ( Xd_0__inst_mult_12_310  ) + ( Xd_0__inst_mult_12_309  ))
// Xd_0__inst_mult_12_433  = CARRY(( (din_a[149] & din_b[144]) ) + ( Xd_0__inst_mult_12_310  ) + ( Xd_0__inst_mult_12_309  ))
// Xd_0__inst_mult_12_434  = SHARE((din_b[144] & din_a[150]))

	.dataa(!din_a[149]),
	.datab(!din_b[144]),
	.datac(!din_a[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_309 ),
	.sharein(Xd_0__inst_mult_12_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_432 ),
	.cout(Xd_0__inst_mult_12_433 ),
	.shareout(Xd_0__inst_mult_12_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_131 (
// Equation(s):
// Xd_0__inst_mult_12_436  = SUM(( (din_a[147] & din_b[146]) ) + ( Xd_0__inst_mult_12_314  ) + ( Xd_0__inst_mult_12_313  ))
// Xd_0__inst_mult_12_437  = CARRY(( (din_a[147] & din_b[146]) ) + ( Xd_0__inst_mult_12_314  ) + ( Xd_0__inst_mult_12_313  ))
// Xd_0__inst_mult_12_438  = SHARE((din_b[146] & din_a[148]))

	.dataa(!din_a[147]),
	.datab(!din_b[146]),
	.datac(!din_a[148]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_313 ),
	.sharein(Xd_0__inst_mult_12_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_436 ),
	.cout(Xd_0__inst_mult_12_437 ),
	.shareout(Xd_0__inst_mult_12_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_59 (
// Equation(s):
// Xd_0__inst_mult_10_59_sumout  = SUM(( (din_a[130] & din_b[120]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_60  = CARRY(( (din_a[130] & din_b[120]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_61  = SHARE(GND)

	.dataa(!din_a[130]),
	.datab(!din_b[120]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_10_59_sumout ),
	.cout(Xd_0__inst_mult_10_60 ),
	.shareout(Xd_0__inst_mult_10_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_127 (
// Equation(s):
// Xd_0__inst_mult_13_408  = SUM(( (din_a[161] & din_b[156]) ) + ( Xd_0__inst_mult_13_290  ) + ( Xd_0__inst_mult_13_289  ))
// Xd_0__inst_mult_13_409  = CARRY(( (din_a[161] & din_b[156]) ) + ( Xd_0__inst_mult_13_290  ) + ( Xd_0__inst_mult_13_289  ))
// Xd_0__inst_mult_13_410  = SHARE((din_b[156] & din_a[162]))

	.dataa(!din_a[161]),
	.datab(!din_b[156]),
	.datac(!din_a[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_289 ),
	.sharein(Xd_0__inst_mult_13_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_408 ),
	.cout(Xd_0__inst_mult_13_409 ),
	.shareout(Xd_0__inst_mult_13_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_128 (
// Equation(s):
// Xd_0__inst_mult_13_412  = SUM(( (din_a[159] & din_b[158]) ) + ( Xd_0__inst_mult_13_294  ) + ( Xd_0__inst_mult_13_293  ))
// Xd_0__inst_mult_13_413  = CARRY(( (din_a[159] & din_b[158]) ) + ( Xd_0__inst_mult_13_294  ) + ( Xd_0__inst_mult_13_293  ))
// Xd_0__inst_mult_13_414  = SHARE((din_b[158] & din_a[160]))

	.dataa(!din_a[159]),
	.datab(!din_b[158]),
	.datac(!din_a[160]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_293 ),
	.sharein(Xd_0__inst_mult_13_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_412 ),
	.cout(Xd_0__inst_mult_13_413 ),
	.shareout(Xd_0__inst_mult_13_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_63 (
// Equation(s):
// Xd_0__inst_mult_15_63_sumout  = SUM(( (din_a[190] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_64  = CARRY(( (din_a[190] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_65  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_15_63_sumout ),
	.cout(Xd_0__inst_mult_15_64 ),
	.shareout(Xd_0__inst_mult_15_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_131 (
// Equation(s):
// Xd_0__inst_mult_14_424  = SUM(( (din_a[173] & din_b[168]) ) + ( Xd_0__inst_mult_14_314  ) + ( Xd_0__inst_mult_14_313  ))
// Xd_0__inst_mult_14_425  = CARRY(( (din_a[173] & din_b[168]) ) + ( Xd_0__inst_mult_14_314  ) + ( Xd_0__inst_mult_14_313  ))
// Xd_0__inst_mult_14_426  = SHARE((din_b[168] & din_a[174]))

	.dataa(!din_a[173]),
	.datab(!din_b[168]),
	.datac(!din_a[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_313 ),
	.sharein(Xd_0__inst_mult_14_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_424 ),
	.cout(Xd_0__inst_mult_14_425 ),
	.shareout(Xd_0__inst_mult_14_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_132 (
// Equation(s):
// Xd_0__inst_mult_14_428  = SUM(( (din_a[171] & din_b[170]) ) + ( Xd_0__inst_mult_14_318  ) + ( Xd_0__inst_mult_14_317  ))
// Xd_0__inst_mult_14_429  = CARRY(( (din_a[171] & din_b[170]) ) + ( Xd_0__inst_mult_14_318  ) + ( Xd_0__inst_mult_14_317  ))
// Xd_0__inst_mult_14_430  = SHARE((din_b[170] & din_a[172]))

	.dataa(!din_a[171]),
	.datab(!din_b[170]),
	.datac(!din_a[172]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_317 ),
	.sharein(Xd_0__inst_mult_14_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_428 ),
	.cout(Xd_0__inst_mult_14_429 ),
	.shareout(Xd_0__inst_mult_14_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_55 (
// Equation(s):
// Xd_0__inst_mult_4_55_sumout  = SUM(( (din_a[58] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_56  = CARRY(( (din_a[58] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_57  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_55_sumout ),
	.cout(Xd_0__inst_mult_4_56 ),
	.shareout(Xd_0__inst_mult_4_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_134 (
// Equation(s):
// Xd_0__inst_mult_15_436  = SUM(( (din_a[185] & din_b[180]) ) + ( Xd_0__inst_mult_15_314  ) + ( Xd_0__inst_mult_15_313  ))
// Xd_0__inst_mult_15_437  = CARRY(( (din_a[185] & din_b[180]) ) + ( Xd_0__inst_mult_15_314  ) + ( Xd_0__inst_mult_15_313  ))
// Xd_0__inst_mult_15_438  = SHARE((din_b[180] & din_a[186]))

	.dataa(!din_a[185]),
	.datab(!din_b[180]),
	.datac(!din_a[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_313 ),
	.sharein(Xd_0__inst_mult_15_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_436 ),
	.cout(Xd_0__inst_mult_15_437 ),
	.shareout(Xd_0__inst_mult_15_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_135 (
// Equation(s):
// Xd_0__inst_mult_15_440  = SUM(( (din_a[183] & din_b[182]) ) + ( Xd_0__inst_mult_15_318  ) + ( Xd_0__inst_mult_15_317  ))
// Xd_0__inst_mult_15_441  = CARRY(( (din_a[183] & din_b[182]) ) + ( Xd_0__inst_mult_15_318  ) + ( Xd_0__inst_mult_15_317  ))
// Xd_0__inst_mult_15_442  = SHARE((din_b[182] & din_a[184]))

	.dataa(!din_a[183]),
	.datab(!din_b[182]),
	.datac(!din_a[184]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_317 ),
	.sharein(Xd_0__inst_mult_15_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_440 ),
	.cout(Xd_0__inst_mult_15_441 ),
	.shareout(Xd_0__inst_mult_15_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_55 (
// Equation(s):
// Xd_0__inst_mult_9_55_sumout  = SUM(( (din_a[118] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_56  = CARRY(( (din_a[118] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_57  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[108]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_55_sumout ),
	.cout(Xd_0__inst_mult_9_56 ),
	.shareout(Xd_0__inst_mult_9_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_123 (
// Equation(s):
// Xd_0__inst_mult_10_404  = SUM(( (din_a[125] & din_b[120]) ) + ( Xd_0__inst_mult_10_286  ) + ( Xd_0__inst_mult_10_285  ))
// Xd_0__inst_mult_10_405  = CARRY(( (din_a[125] & din_b[120]) ) + ( Xd_0__inst_mult_10_286  ) + ( Xd_0__inst_mult_10_285  ))
// Xd_0__inst_mult_10_406  = SHARE((din_b[120] & din_a[126]))

	.dataa(!din_a[125]),
	.datab(!din_b[120]),
	.datac(!din_a[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_285 ),
	.sharein(Xd_0__inst_mult_10_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_404 ),
	.cout(Xd_0__inst_mult_10_405 ),
	.shareout(Xd_0__inst_mult_10_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_124 (
// Equation(s):
// Xd_0__inst_mult_10_408  = SUM(( (din_a[123] & din_b[122]) ) + ( Xd_0__inst_mult_10_290  ) + ( Xd_0__inst_mult_10_289  ))
// Xd_0__inst_mult_10_409  = CARRY(( (din_a[123] & din_b[122]) ) + ( Xd_0__inst_mult_10_290  ) + ( Xd_0__inst_mult_10_289  ))
// Xd_0__inst_mult_10_410  = SHARE((din_b[122] & din_a[124]))

	.dataa(!din_a[123]),
	.datab(!din_b[122]),
	.datac(!din_a[124]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_289 ),
	.sharein(Xd_0__inst_mult_10_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_408 ),
	.cout(Xd_0__inst_mult_10_409 ),
	.shareout(Xd_0__inst_mult_10_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_59 (
// Equation(s):
// Xd_0__inst_mult_0_59_sumout  = SUM(( (din_a[9] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_60  = CARRY(( (din_a[9] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_61  = SHARE(GND)

	.dataa(!din_a[9]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_59_sumout ),
	.cout(Xd_0__inst_mult_0_60 ),
	.shareout(Xd_0__inst_mult_0_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_127 (
// Equation(s):
// Xd_0__inst_mult_11_408  = SUM(( (din_a[137] & din_b[132]) ) + ( Xd_0__inst_mult_11_290  ) + ( Xd_0__inst_mult_11_289  ))
// Xd_0__inst_mult_11_409  = CARRY(( (din_a[137] & din_b[132]) ) + ( Xd_0__inst_mult_11_290  ) + ( Xd_0__inst_mult_11_289  ))
// Xd_0__inst_mult_11_410  = SHARE((din_b[132] & din_a[138]))

	.dataa(!din_a[137]),
	.datab(!din_b[132]),
	.datac(!din_a[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_289 ),
	.sharein(Xd_0__inst_mult_11_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_408 ),
	.cout(Xd_0__inst_mult_11_409 ),
	.shareout(Xd_0__inst_mult_11_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_128 (
// Equation(s):
// Xd_0__inst_mult_11_412  = SUM(( (din_a[135] & din_b[134]) ) + ( Xd_0__inst_mult_11_294  ) + ( Xd_0__inst_mult_11_293  ))
// Xd_0__inst_mult_11_413  = CARRY(( (din_a[135] & din_b[134]) ) + ( Xd_0__inst_mult_11_294  ) + ( Xd_0__inst_mult_11_293  ))
// Xd_0__inst_mult_11_414  = SHARE((din_b[134] & din_a[136]))

	.dataa(!din_a[135]),
	.datab(!din_b[134]),
	.datac(!din_a[136]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_293 ),
	.sharein(Xd_0__inst_mult_11_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_412 ),
	.cout(Xd_0__inst_mult_11_413 ),
	.shareout(Xd_0__inst_mult_11_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_55 (
// Equation(s):
// Xd_0__inst_mult_11_55_sumout  = SUM(( (din_a[142] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_56  = CARRY(( (din_a[142] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_57  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_55_sumout ),
	.cout(Xd_0__inst_mult_11_56 ),
	.shareout(Xd_0__inst_mult_11_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_127 (
// Equation(s):
// Xd_0__inst_mult_8_408  = SUM(( (din_a[101] & din_b[96]) ) + ( Xd_0__inst_mult_8_290  ) + ( Xd_0__inst_mult_8_289  ))
// Xd_0__inst_mult_8_409  = CARRY(( (din_a[101] & din_b[96]) ) + ( Xd_0__inst_mult_8_290  ) + ( Xd_0__inst_mult_8_289  ))
// Xd_0__inst_mult_8_410  = SHARE((din_b[96] & din_a[102]))

	.dataa(!din_a[101]),
	.datab(!din_b[96]),
	.datac(!din_a[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_289 ),
	.sharein(Xd_0__inst_mult_8_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_408 ),
	.cout(Xd_0__inst_mult_8_409 ),
	.shareout(Xd_0__inst_mult_8_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_128 (
// Equation(s):
// Xd_0__inst_mult_8_412  = SUM(( (din_a[99] & din_b[98]) ) + ( Xd_0__inst_mult_8_294  ) + ( Xd_0__inst_mult_8_293  ))
// Xd_0__inst_mult_8_413  = CARRY(( (din_a[99] & din_b[98]) ) + ( Xd_0__inst_mult_8_294  ) + ( Xd_0__inst_mult_8_293  ))
// Xd_0__inst_mult_8_414  = SHARE((din_b[98] & din_a[100]))

	.dataa(!din_a[99]),
	.datab(!din_b[98]),
	.datac(!din_a[100]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_293 ),
	.sharein(Xd_0__inst_mult_8_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_412 ),
	.cout(Xd_0__inst_mult_8_413 ),
	.shareout(Xd_0__inst_mult_8_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_123 (
// Equation(s):
// Xd_0__inst_mult_9_404  = SUM(( (din_a[113] & din_b[108]) ) + ( Xd_0__inst_mult_9_286  ) + ( Xd_0__inst_mult_9_285  ))
// Xd_0__inst_mult_9_405  = CARRY(( (din_a[113] & din_b[108]) ) + ( Xd_0__inst_mult_9_286  ) + ( Xd_0__inst_mult_9_285  ))
// Xd_0__inst_mult_9_406  = SHARE((din_b[108] & din_a[114]))

	.dataa(!din_a[113]),
	.datab(!din_b[108]),
	.datac(!din_a[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_285 ),
	.sharein(Xd_0__inst_mult_9_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_404 ),
	.cout(Xd_0__inst_mult_9_405 ),
	.shareout(Xd_0__inst_mult_9_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_124 (
// Equation(s):
// Xd_0__inst_mult_9_408  = SUM(( (din_a[111] & din_b[110]) ) + ( Xd_0__inst_mult_9_290  ) + ( Xd_0__inst_mult_9_289  ))
// Xd_0__inst_mult_9_409  = CARRY(( (din_a[111] & din_b[110]) ) + ( Xd_0__inst_mult_9_290  ) + ( Xd_0__inst_mult_9_289  ))
// Xd_0__inst_mult_9_410  = SHARE((din_b[110] & din_a[112]))

	.dataa(!din_a[111]),
	.datab(!din_b[110]),
	.datac(!din_a[112]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_289 ),
	.sharein(Xd_0__inst_mult_9_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_408 ),
	.cout(Xd_0__inst_mult_9_409 ),
	.shareout(Xd_0__inst_mult_9_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_123 (
// Equation(s):
// Xd_0__inst_mult_6_404  = SUM(( (din_a[77] & din_b[72]) ) + ( Xd_0__inst_mult_6_286  ) + ( Xd_0__inst_mult_6_285  ))
// Xd_0__inst_mult_6_405  = CARRY(( (din_a[77] & din_b[72]) ) + ( Xd_0__inst_mult_6_286  ) + ( Xd_0__inst_mult_6_285  ))
// Xd_0__inst_mult_6_406  = SHARE((din_b[72] & din_a[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[72]),
	.datac(!din_a[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_285 ),
	.sharein(Xd_0__inst_mult_6_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_404 ),
	.cout(Xd_0__inst_mult_6_405 ),
	.shareout(Xd_0__inst_mult_6_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_124 (
// Equation(s):
// Xd_0__inst_mult_6_408  = SUM(( (din_a[75] & din_b[74]) ) + ( Xd_0__inst_mult_6_290  ) + ( Xd_0__inst_mult_6_289  ))
// Xd_0__inst_mult_6_409  = CARRY(( (din_a[75] & din_b[74]) ) + ( Xd_0__inst_mult_6_290  ) + ( Xd_0__inst_mult_6_289  ))
// Xd_0__inst_mult_6_410  = SHARE((din_b[74] & din_a[76]))

	.dataa(!din_a[75]),
	.datab(!din_b[74]),
	.datac(!din_a[76]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_289 ),
	.sharein(Xd_0__inst_mult_6_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_408 ),
	.cout(Xd_0__inst_mult_6_409 ),
	.shareout(Xd_0__inst_mult_6_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_119 (
// Equation(s):
// Xd_0__inst_mult_7_388  = SUM(( (din_a[89] & din_b[84]) ) + ( Xd_0__inst_mult_7_262  ) + ( Xd_0__inst_mult_7_261  ))
// Xd_0__inst_mult_7_389  = CARRY(( (din_a[89] & din_b[84]) ) + ( Xd_0__inst_mult_7_262  ) + ( Xd_0__inst_mult_7_261  ))
// Xd_0__inst_mult_7_390  = SHARE((din_b[84] & din_a[90]))

	.dataa(!din_a[89]),
	.datab(!din_b[84]),
	.datac(!din_a[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_261 ),
	.sharein(Xd_0__inst_mult_7_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_388 ),
	.cout(Xd_0__inst_mult_7_389 ),
	.shareout(Xd_0__inst_mult_7_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_120 (
// Equation(s):
// Xd_0__inst_mult_7_392  = SUM(( (din_a[87] & din_b[86]) ) + ( Xd_0__inst_mult_7_266  ) + ( Xd_0__inst_mult_7_265  ))
// Xd_0__inst_mult_7_393  = CARRY(( (din_a[87] & din_b[86]) ) + ( Xd_0__inst_mult_7_266  ) + ( Xd_0__inst_mult_7_265  ))
// Xd_0__inst_mult_7_394  = SHARE((din_b[86] & din_a[88]))

	.dataa(!din_a[87]),
	.datab(!din_b[86]),
	.datac(!din_a[88]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_265 ),
	.sharein(Xd_0__inst_mult_7_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_392 ),
	.cout(Xd_0__inst_mult_7_393 ),
	.shareout(Xd_0__inst_mult_7_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_132 (
// Equation(s):
// Xd_0__inst_mult_4_428  = SUM(( (din_a[53] & din_b[48]) ) + ( Xd_0__inst_mult_4_298  ) + ( Xd_0__inst_mult_4_297  ))
// Xd_0__inst_mult_4_429  = CARRY(( (din_a[53] & din_b[48]) ) + ( Xd_0__inst_mult_4_298  ) + ( Xd_0__inst_mult_4_297  ))
// Xd_0__inst_mult_4_430  = SHARE((din_b[48] & din_a[54]))

	.dataa(!din_a[53]),
	.datab(!din_b[48]),
	.datac(!din_a[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_297 ),
	.sharein(Xd_0__inst_mult_4_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_428 ),
	.cout(Xd_0__inst_mult_4_429 ),
	.shareout(Xd_0__inst_mult_4_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_133 (
// Equation(s):
// Xd_0__inst_mult_4_432  = SUM(( (din_a[51] & din_b[50]) ) + ( Xd_0__inst_mult_4_302  ) + ( Xd_0__inst_mult_4_301  ))
// Xd_0__inst_mult_4_433  = CARRY(( (din_a[51] & din_b[50]) ) + ( Xd_0__inst_mult_4_302  ) + ( Xd_0__inst_mult_4_301  ))
// Xd_0__inst_mult_4_434  = SHARE((din_b[50] & din_a[52]))

	.dataa(!din_a[51]),
	.datab(!din_b[50]),
	.datac(!din_a[52]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_301 ),
	.sharein(Xd_0__inst_mult_4_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_432 ),
	.cout(Xd_0__inst_mult_4_433 ),
	.shareout(Xd_0__inst_mult_4_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_59 (
// Equation(s):
// Xd_0__inst_mult_2_59_sumout  = SUM(( (din_a[31] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_60  = CARRY(( (din_a[31] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_61  = SHARE(GND)

	.dataa(!din_a[31]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_59_sumout ),
	.cout(Xd_0__inst_mult_2_60 ),
	.shareout(Xd_0__inst_mult_2_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_119 (
// Equation(s):
// Xd_0__inst_mult_5_388  = SUM(( (din_a[65] & din_b[60]) ) + ( Xd_0__inst_mult_5_262  ) + ( Xd_0__inst_mult_5_261  ))
// Xd_0__inst_mult_5_389  = CARRY(( (din_a[65] & din_b[60]) ) + ( Xd_0__inst_mult_5_262  ) + ( Xd_0__inst_mult_5_261  ))
// Xd_0__inst_mult_5_390  = SHARE((din_b[60] & din_a[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[60]),
	.datac(!din_a[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_261 ),
	.sharein(Xd_0__inst_mult_5_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_388 ),
	.cout(Xd_0__inst_mult_5_389 ),
	.shareout(Xd_0__inst_mult_5_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_120 (
// Equation(s):
// Xd_0__inst_mult_5_392  = SUM(( (din_a[63] & din_b[62]) ) + ( Xd_0__inst_mult_5_266  ) + ( Xd_0__inst_mult_5_265  ))
// Xd_0__inst_mult_5_393  = CARRY(( (din_a[63] & din_b[62]) ) + ( Xd_0__inst_mult_5_266  ) + ( Xd_0__inst_mult_5_265  ))
// Xd_0__inst_mult_5_394  = SHARE((din_b[62] & din_a[64]))

	.dataa(!din_a[63]),
	.datab(!din_b[62]),
	.datac(!din_a[64]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_265 ),
	.sharein(Xd_0__inst_mult_5_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_392 ),
	.cout(Xd_0__inst_mult_5_393 ),
	.shareout(Xd_0__inst_mult_5_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_123 (
// Equation(s):
// Xd_0__inst_mult_2_392  = SUM(( (din_a[29] & din_b[24]) ) + ( Xd_0__inst_mult_2_266  ) + ( Xd_0__inst_mult_2_265  ))
// Xd_0__inst_mult_2_393  = CARRY(( (din_a[29] & din_b[24]) ) + ( Xd_0__inst_mult_2_266  ) + ( Xd_0__inst_mult_2_265  ))
// Xd_0__inst_mult_2_394  = SHARE((din_b[24] & din_a[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[24]),
	.datac(!din_a[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_265 ),
	.sharein(Xd_0__inst_mult_2_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_392 ),
	.cout(Xd_0__inst_mult_2_393 ),
	.shareout(Xd_0__inst_mult_2_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_124 (
// Equation(s):
// Xd_0__inst_mult_2_396  = SUM(( (din_a[27] & din_b[26]) ) + ( Xd_0__inst_mult_2_270  ) + ( Xd_0__inst_mult_2_269  ))
// Xd_0__inst_mult_2_397  = CARRY(( (din_a[27] & din_b[26]) ) + ( Xd_0__inst_mult_2_270  ) + ( Xd_0__inst_mult_2_269  ))
// Xd_0__inst_mult_2_398  = SHARE((din_b[26] & din_a[28]))

	.dataa(!din_a[27]),
	.datab(!din_b[26]),
	.datac(!din_a[28]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_269 ),
	.sharein(Xd_0__inst_mult_2_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_396 ),
	.cout(Xd_0__inst_mult_2_397 ),
	.shareout(Xd_0__inst_mult_2_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_119 (
// Equation(s):
// Xd_0__inst_mult_3_388  = SUM(( (din_a[41] & din_b[36]) ) + ( Xd_0__inst_mult_3_262  ) + ( Xd_0__inst_mult_3_261  ))
// Xd_0__inst_mult_3_389  = CARRY(( (din_a[41] & din_b[36]) ) + ( Xd_0__inst_mult_3_262  ) + ( Xd_0__inst_mult_3_261  ))
// Xd_0__inst_mult_3_390  = SHARE((din_b[36] & din_a[42]))

	.dataa(!din_a[41]),
	.datab(!din_b[36]),
	.datac(!din_a[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_261 ),
	.sharein(Xd_0__inst_mult_3_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_388 ),
	.cout(Xd_0__inst_mult_3_389 ),
	.shareout(Xd_0__inst_mult_3_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_120 (
// Equation(s):
// Xd_0__inst_mult_3_392  = SUM(( (din_a[39] & din_b[38]) ) + ( Xd_0__inst_mult_3_266  ) + ( Xd_0__inst_mult_3_265  ))
// Xd_0__inst_mult_3_393  = CARRY(( (din_a[39] & din_b[38]) ) + ( Xd_0__inst_mult_3_266  ) + ( Xd_0__inst_mult_3_265  ))
// Xd_0__inst_mult_3_394  = SHARE((din_b[38] & din_a[40]))

	.dataa(!din_a[39]),
	.datab(!din_b[38]),
	.datac(!din_a[40]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_265 ),
	.sharein(Xd_0__inst_mult_3_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_392 ),
	.cout(Xd_0__inst_mult_3_393 ),
	.shareout(Xd_0__inst_mult_3_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_59 (
// Equation(s):
// Xd_0__inst_mult_11_59_sumout  = SUM(( (din_a[140] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_60  = CARRY(( (din_a[140] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_61  = SHARE(GND)

	.dataa(!din_a[140]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_59_sumout ),
	.cout(Xd_0__inst_mult_11_60 ),
	.shareout(Xd_0__inst_mult_11_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_123 (
// Equation(s):
// Xd_0__inst_mult_0_392  = SUM(( (din_a[5] & din_b[0]) ) + ( Xd_0__inst_mult_0_266  ) + ( Xd_0__inst_mult_0_265  ))
// Xd_0__inst_mult_0_393  = CARRY(( (din_a[5] & din_b[0]) ) + ( Xd_0__inst_mult_0_266  ) + ( Xd_0__inst_mult_0_265  ))
// Xd_0__inst_mult_0_394  = SHARE((din_b[0] & din_a[6]))

	.dataa(!din_a[5]),
	.datab(!din_b[0]),
	.datac(!din_a[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_265 ),
	.sharein(Xd_0__inst_mult_0_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_392 ),
	.cout(Xd_0__inst_mult_0_393 ),
	.shareout(Xd_0__inst_mult_0_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_124 (
// Equation(s):
// Xd_0__inst_mult_0_396  = SUM(( (din_a[3] & din_b[2]) ) + ( Xd_0__inst_mult_0_270  ) + ( Xd_0__inst_mult_0_269  ))
// Xd_0__inst_mult_0_397  = CARRY(( (din_a[3] & din_b[2]) ) + ( Xd_0__inst_mult_0_270  ) + ( Xd_0__inst_mult_0_269  ))
// Xd_0__inst_mult_0_398  = SHARE((din_b[2] & din_a[4]))

	.dataa(!din_a[3]),
	.datab(!din_b[2]),
	.datac(!din_a[4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_269 ),
	.sharein(Xd_0__inst_mult_0_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_396 ),
	.cout(Xd_0__inst_mult_0_397 ),
	.shareout(Xd_0__inst_mult_0_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_63 (
// Equation(s):
// Xd_0__inst_mult_12_63_sumout  = SUM(( (din_a[152] & din_b[144]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_64  = CARRY(( (din_a[152] & din_b[144]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_65  = SHARE(GND)

	.dataa(!din_a[152]),
	.datab(!din_b[144]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_12_63_sumout ),
	.cout(Xd_0__inst_mult_12_64 ),
	.shareout(Xd_0__inst_mult_12_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_123 (
// Equation(s):
// Xd_0__inst_mult_1_392  = SUM(( (din_a[17] & din_b[12]) ) + ( Xd_0__inst_mult_1_266  ) + ( Xd_0__inst_mult_1_265  ))
// Xd_0__inst_mult_1_393  = CARRY(( (din_a[17] & din_b[12]) ) + ( Xd_0__inst_mult_1_266  ) + ( Xd_0__inst_mult_1_265  ))
// Xd_0__inst_mult_1_394  = SHARE((din_b[12] & din_a[18]))

	.dataa(!din_a[17]),
	.datab(!din_b[12]),
	.datac(!din_a[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_265 ),
	.sharein(Xd_0__inst_mult_1_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_392 ),
	.cout(Xd_0__inst_mult_1_393 ),
	.shareout(Xd_0__inst_mult_1_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_124 (
// Equation(s):
// Xd_0__inst_mult_1_396  = SUM(( (din_a[15] & din_b[14]) ) + ( Xd_0__inst_mult_1_270  ) + ( Xd_0__inst_mult_1_269  ))
// Xd_0__inst_mult_1_397  = CARRY(( (din_a[15] & din_b[14]) ) + ( Xd_0__inst_mult_1_270  ) + ( Xd_0__inst_mult_1_269  ))
// Xd_0__inst_mult_1_398  = SHARE((din_b[14] & din_a[16]))

	.dataa(!din_a[15]),
	.datab(!din_b[14]),
	.datac(!din_a[16]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_269 ),
	.sharein(Xd_0__inst_mult_1_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_396 ),
	.cout(Xd_0__inst_mult_1_397 ),
	.shareout(Xd_0__inst_mult_1_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_63 (
// Equation(s):
// Xd_0__inst_mult_1_63_sumout  = SUM(( (din_a[19] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_64  = CARRY(( (din_a[19] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_65  = SHARE(GND)

	.dataa(!din_a[19]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_63_sumout ),
	.cout(Xd_0__inst_mult_1_64 ),
	.shareout(Xd_0__inst_mult_1_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_132 (
// Equation(s):
// Xd_0__inst_mult_12_440  = SUM(( (din_a[149] & din_b[145]) ) + ( Xd_0__inst_mult_12_434  ) + ( Xd_0__inst_mult_12_433  ))
// Xd_0__inst_mult_12_441  = CARRY(( (din_a[149] & din_b[145]) ) + ( Xd_0__inst_mult_12_434  ) + ( Xd_0__inst_mult_12_433  ))
// Xd_0__inst_mult_12_442  = SHARE((din_b[145] & din_a[150]))

	.dataa(!din_a[149]),
	.datab(!din_b[145]),
	.datac(!din_a[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_433 ),
	.sharein(Xd_0__inst_mult_12_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_440 ),
	.cout(Xd_0__inst_mult_12_441 ),
	.shareout(Xd_0__inst_mult_12_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_133 (
// Equation(s):
// Xd_0__inst_mult_12_444  = SUM(( (!din_a[147] & (((din_a[146] & din_b[148])))) # (din_a[147] & (!din_b[147] $ (((!din_a[146]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_438  ) + ( Xd_0__inst_mult_12_437  ))
// Xd_0__inst_mult_12_445  = CARRY(( (!din_a[147] & (((din_a[146] & din_b[148])))) # (din_a[147] & (!din_b[147] $ (((!din_a[146]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_438  ) + ( Xd_0__inst_mult_12_437  ))
// Xd_0__inst_mult_12_446  = SHARE((din_a[147] & (din_b[147] & (din_a[146] & din_b[148]))))

	.dataa(!din_a[147]),
	.datab(!din_b[147]),
	.datac(!din_a[146]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_437 ),
	.sharein(Xd_0__inst_mult_12_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_444 ),
	.cout(Xd_0__inst_mult_12_445 ),
	.shareout(Xd_0__inst_mult_12_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_129 (
// Equation(s):
// Xd_0__inst_mult_13_416  = SUM(( (din_a[161] & din_b[157]) ) + ( Xd_0__inst_mult_13_410  ) + ( Xd_0__inst_mult_13_409  ))
// Xd_0__inst_mult_13_417  = CARRY(( (din_a[161] & din_b[157]) ) + ( Xd_0__inst_mult_13_410  ) + ( Xd_0__inst_mult_13_409  ))
// Xd_0__inst_mult_13_418  = SHARE((din_b[157] & din_a[162]))

	.dataa(!din_a[161]),
	.datab(!din_b[157]),
	.datac(!din_a[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_409 ),
	.sharein(Xd_0__inst_mult_13_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_416 ),
	.cout(Xd_0__inst_mult_13_417 ),
	.shareout(Xd_0__inst_mult_13_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_130 (
// Equation(s):
// Xd_0__inst_mult_13_420  = SUM(( (!din_a[159] & (((din_a[158] & din_b[160])))) # (din_a[159] & (!din_b[159] $ (((!din_a[158]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_414  ) + ( Xd_0__inst_mult_13_413  ))
// Xd_0__inst_mult_13_421  = CARRY(( (!din_a[159] & (((din_a[158] & din_b[160])))) # (din_a[159] & (!din_b[159] $ (((!din_a[158]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_414  ) + ( Xd_0__inst_mult_13_413  ))
// Xd_0__inst_mult_13_422  = SHARE((din_a[159] & (din_b[159] & (din_a[158] & din_b[160]))))

	.dataa(!din_a[159]),
	.datab(!din_b[159]),
	.datac(!din_a[158]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_413 ),
	.sharein(Xd_0__inst_mult_13_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_420 ),
	.cout(Xd_0__inst_mult_13_421 ),
	.shareout(Xd_0__inst_mult_13_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_133 (
// Equation(s):
// Xd_0__inst_mult_14_432  = SUM(( (din_a[173] & din_b[169]) ) + ( Xd_0__inst_mult_14_426  ) + ( Xd_0__inst_mult_14_425  ))
// Xd_0__inst_mult_14_433  = CARRY(( (din_a[173] & din_b[169]) ) + ( Xd_0__inst_mult_14_426  ) + ( Xd_0__inst_mult_14_425  ))
// Xd_0__inst_mult_14_434  = SHARE((din_b[169] & din_a[174]))

	.dataa(!din_a[173]),
	.datab(!din_b[169]),
	.datac(!din_a[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_425 ),
	.sharein(Xd_0__inst_mult_14_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_432 ),
	.cout(Xd_0__inst_mult_14_433 ),
	.shareout(Xd_0__inst_mult_14_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_134 (
// Equation(s):
// Xd_0__inst_mult_14_436  = SUM(( (!din_a[171] & (((din_a[170] & din_b[172])))) # (din_a[171] & (!din_b[171] $ (((!din_a[170]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_430  ) + ( Xd_0__inst_mult_14_429  ))
// Xd_0__inst_mult_14_437  = CARRY(( (!din_a[171] & (((din_a[170] & din_b[172])))) # (din_a[171] & (!din_b[171] $ (((!din_a[170]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_430  ) + ( Xd_0__inst_mult_14_429  ))
// Xd_0__inst_mult_14_438  = SHARE((din_a[171] & (din_b[171] & (din_a[170] & din_b[172]))))

	.dataa(!din_a[171]),
	.datab(!din_b[171]),
	.datac(!din_a[170]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_429 ),
	.sharein(Xd_0__inst_mult_14_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_436 ),
	.cout(Xd_0__inst_mult_14_437 ),
	.shareout(Xd_0__inst_mult_14_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_136 (
// Equation(s):
// Xd_0__inst_mult_15_444  = SUM(( (din_a[185] & din_b[181]) ) + ( Xd_0__inst_mult_15_438  ) + ( Xd_0__inst_mult_15_437  ))
// Xd_0__inst_mult_15_445  = CARRY(( (din_a[185] & din_b[181]) ) + ( Xd_0__inst_mult_15_438  ) + ( Xd_0__inst_mult_15_437  ))
// Xd_0__inst_mult_15_446  = SHARE((din_b[181] & din_a[186]))

	.dataa(!din_a[185]),
	.datab(!din_b[181]),
	.datac(!din_a[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_437 ),
	.sharein(Xd_0__inst_mult_15_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_444 ),
	.cout(Xd_0__inst_mult_15_445 ),
	.shareout(Xd_0__inst_mult_15_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_137 (
// Equation(s):
// Xd_0__inst_mult_15_448  = SUM(( (!din_a[183] & (((din_a[182] & din_b[184])))) # (din_a[183] & (!din_b[183] $ (((!din_a[182]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_442  ) + ( Xd_0__inst_mult_15_441  ))
// Xd_0__inst_mult_15_449  = CARRY(( (!din_a[183] & (((din_a[182] & din_b[184])))) # (din_a[183] & (!din_b[183] $ (((!din_a[182]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_442  ) + ( Xd_0__inst_mult_15_441  ))
// Xd_0__inst_mult_15_450  = SHARE((din_a[183] & (din_b[183] & (din_a[182] & din_b[184]))))

	.dataa(!din_a[183]),
	.datab(!din_b[183]),
	.datac(!din_a[182]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_441 ),
	.sharein(Xd_0__inst_mult_15_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_448 ),
	.cout(Xd_0__inst_mult_15_449 ),
	.shareout(Xd_0__inst_mult_15_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_125 (
// Equation(s):
// Xd_0__inst_mult_10_412  = SUM(( (din_a[125] & din_b[121]) ) + ( Xd_0__inst_mult_10_406  ) + ( Xd_0__inst_mult_10_405  ))
// Xd_0__inst_mult_10_413  = CARRY(( (din_a[125] & din_b[121]) ) + ( Xd_0__inst_mult_10_406  ) + ( Xd_0__inst_mult_10_405  ))
// Xd_0__inst_mult_10_414  = SHARE((din_b[121] & din_a[126]))

	.dataa(!din_a[125]),
	.datab(!din_b[121]),
	.datac(!din_a[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_405 ),
	.sharein(Xd_0__inst_mult_10_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_412 ),
	.cout(Xd_0__inst_mult_10_413 ),
	.shareout(Xd_0__inst_mult_10_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_126 (
// Equation(s):
// Xd_0__inst_mult_10_416  = SUM(( (!din_a[123] & (((din_a[122] & din_b[124])))) # (din_a[123] & (!din_b[123] $ (((!din_a[122]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_410  ) + ( Xd_0__inst_mult_10_409  ))
// Xd_0__inst_mult_10_417  = CARRY(( (!din_a[123] & (((din_a[122] & din_b[124])))) # (din_a[123] & (!din_b[123] $ (((!din_a[122]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_410  ) + ( Xd_0__inst_mult_10_409  ))
// Xd_0__inst_mult_10_418  = SHARE((din_a[123] & (din_b[123] & (din_a[122] & din_b[124]))))

	.dataa(!din_a[123]),
	.datab(!din_b[123]),
	.datac(!din_a[122]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_409 ),
	.sharein(Xd_0__inst_mult_10_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_416 ),
	.cout(Xd_0__inst_mult_10_417 ),
	.shareout(Xd_0__inst_mult_10_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_129 (
// Equation(s):
// Xd_0__inst_mult_11_416  = SUM(( (din_a[137] & din_b[133]) ) + ( Xd_0__inst_mult_11_410  ) + ( Xd_0__inst_mult_11_409  ))
// Xd_0__inst_mult_11_417  = CARRY(( (din_a[137] & din_b[133]) ) + ( Xd_0__inst_mult_11_410  ) + ( Xd_0__inst_mult_11_409  ))
// Xd_0__inst_mult_11_418  = SHARE((din_b[133] & din_a[138]))

	.dataa(!din_a[137]),
	.datab(!din_b[133]),
	.datac(!din_a[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_409 ),
	.sharein(Xd_0__inst_mult_11_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_416 ),
	.cout(Xd_0__inst_mult_11_417 ),
	.shareout(Xd_0__inst_mult_11_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_130 (
// Equation(s):
// Xd_0__inst_mult_11_420  = SUM(( (!din_a[135] & (((din_a[134] & din_b[136])))) # (din_a[135] & (!din_b[135] $ (((!din_a[134]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_414  ) + ( Xd_0__inst_mult_11_413  ))
// Xd_0__inst_mult_11_421  = CARRY(( (!din_a[135] & (((din_a[134] & din_b[136])))) # (din_a[135] & (!din_b[135] $ (((!din_a[134]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_414  ) + ( Xd_0__inst_mult_11_413  ))
// Xd_0__inst_mult_11_422  = SHARE((din_a[135] & (din_b[135] & (din_a[134] & din_b[136]))))

	.dataa(!din_a[135]),
	.datab(!din_b[135]),
	.datac(!din_a[134]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_413 ),
	.sharein(Xd_0__inst_mult_11_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_420 ),
	.cout(Xd_0__inst_mult_11_421 ),
	.shareout(Xd_0__inst_mult_11_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_129 (
// Equation(s):
// Xd_0__inst_mult_8_416  = SUM(( (din_a[101] & din_b[97]) ) + ( Xd_0__inst_mult_8_410  ) + ( Xd_0__inst_mult_8_409  ))
// Xd_0__inst_mult_8_417  = CARRY(( (din_a[101] & din_b[97]) ) + ( Xd_0__inst_mult_8_410  ) + ( Xd_0__inst_mult_8_409  ))
// Xd_0__inst_mult_8_418  = SHARE((din_b[97] & din_a[102]))

	.dataa(!din_a[101]),
	.datab(!din_b[97]),
	.datac(!din_a[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_409 ),
	.sharein(Xd_0__inst_mult_8_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_416 ),
	.cout(Xd_0__inst_mult_8_417 ),
	.shareout(Xd_0__inst_mult_8_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_130 (
// Equation(s):
// Xd_0__inst_mult_8_420  = SUM(( (!din_a[99] & (((din_a[98] & din_b[100])))) # (din_a[99] & (!din_b[99] $ (((!din_a[98]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_414  ) + ( Xd_0__inst_mult_8_413  ))
// Xd_0__inst_mult_8_421  = CARRY(( (!din_a[99] & (((din_a[98] & din_b[100])))) # (din_a[99] & (!din_b[99] $ (((!din_a[98]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_414  ) + ( Xd_0__inst_mult_8_413  ))
// Xd_0__inst_mult_8_422  = SHARE((din_a[99] & (din_b[99] & (din_a[98] & din_b[100]))))

	.dataa(!din_a[99]),
	.datab(!din_b[99]),
	.datac(!din_a[98]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_413 ),
	.sharein(Xd_0__inst_mult_8_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_420 ),
	.cout(Xd_0__inst_mult_8_421 ),
	.shareout(Xd_0__inst_mult_8_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_125 (
// Equation(s):
// Xd_0__inst_mult_9_412  = SUM(( (din_a[113] & din_b[109]) ) + ( Xd_0__inst_mult_9_406  ) + ( Xd_0__inst_mult_9_405  ))
// Xd_0__inst_mult_9_413  = CARRY(( (din_a[113] & din_b[109]) ) + ( Xd_0__inst_mult_9_406  ) + ( Xd_0__inst_mult_9_405  ))
// Xd_0__inst_mult_9_414  = SHARE((din_b[109] & din_a[114]))

	.dataa(!din_a[113]),
	.datab(!din_b[109]),
	.datac(!din_a[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_405 ),
	.sharein(Xd_0__inst_mult_9_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_412 ),
	.cout(Xd_0__inst_mult_9_413 ),
	.shareout(Xd_0__inst_mult_9_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_126 (
// Equation(s):
// Xd_0__inst_mult_9_416  = SUM(( (!din_a[111] & (((din_a[110] & din_b[112])))) # (din_a[111] & (!din_b[111] $ (((!din_a[110]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_410  ) + ( Xd_0__inst_mult_9_409  ))
// Xd_0__inst_mult_9_417  = CARRY(( (!din_a[111] & (((din_a[110] & din_b[112])))) # (din_a[111] & (!din_b[111] $ (((!din_a[110]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_410  ) + ( Xd_0__inst_mult_9_409  ))
// Xd_0__inst_mult_9_418  = SHARE((din_a[111] & (din_b[111] & (din_a[110] & din_b[112]))))

	.dataa(!din_a[111]),
	.datab(!din_b[111]),
	.datac(!din_a[110]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_409 ),
	.sharein(Xd_0__inst_mult_9_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_416 ),
	.cout(Xd_0__inst_mult_9_417 ),
	.shareout(Xd_0__inst_mult_9_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_125 (
// Equation(s):
// Xd_0__inst_mult_6_412  = SUM(( (din_a[77] & din_b[73]) ) + ( Xd_0__inst_mult_6_406  ) + ( Xd_0__inst_mult_6_405  ))
// Xd_0__inst_mult_6_413  = CARRY(( (din_a[77] & din_b[73]) ) + ( Xd_0__inst_mult_6_406  ) + ( Xd_0__inst_mult_6_405  ))
// Xd_0__inst_mult_6_414  = SHARE((din_b[73] & din_a[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[73]),
	.datac(!din_a[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_405 ),
	.sharein(Xd_0__inst_mult_6_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_412 ),
	.cout(Xd_0__inst_mult_6_413 ),
	.shareout(Xd_0__inst_mult_6_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_126 (
// Equation(s):
// Xd_0__inst_mult_6_416  = SUM(( (!din_a[75] & (((din_a[74] & din_b[76])))) # (din_a[75] & (!din_b[75] $ (((!din_a[74]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_410  ) + ( Xd_0__inst_mult_6_409  ))
// Xd_0__inst_mult_6_417  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[76])))) # (din_a[75] & (!din_b[75] $ (((!din_a[74]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_410  ) + ( Xd_0__inst_mult_6_409  ))
// Xd_0__inst_mult_6_418  = SHARE((din_a[75] & (din_b[75] & (din_a[74] & din_b[76]))))

	.dataa(!din_a[75]),
	.datab(!din_b[75]),
	.datac(!din_a[74]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_409 ),
	.sharein(Xd_0__inst_mult_6_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_416 ),
	.cout(Xd_0__inst_mult_6_417 ),
	.shareout(Xd_0__inst_mult_6_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_121 (
// Equation(s):
// Xd_0__inst_mult_7_396  = SUM(( (din_a[89] & din_b[85]) ) + ( Xd_0__inst_mult_7_390  ) + ( Xd_0__inst_mult_7_389  ))
// Xd_0__inst_mult_7_397  = CARRY(( (din_a[89] & din_b[85]) ) + ( Xd_0__inst_mult_7_390  ) + ( Xd_0__inst_mult_7_389  ))
// Xd_0__inst_mult_7_398  = SHARE((din_b[85] & din_a[90]))

	.dataa(!din_a[89]),
	.datab(!din_b[85]),
	.datac(!din_a[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_389 ),
	.sharein(Xd_0__inst_mult_7_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_396 ),
	.cout(Xd_0__inst_mult_7_397 ),
	.shareout(Xd_0__inst_mult_7_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_122 (
// Equation(s):
// Xd_0__inst_mult_7_400  = SUM(( (!din_a[87] & (((din_a[86] & din_b[88])))) # (din_a[87] & (!din_b[87] $ (((!din_a[86]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_394  ) + ( Xd_0__inst_mult_7_393  ))
// Xd_0__inst_mult_7_401  = CARRY(( (!din_a[87] & (((din_a[86] & din_b[88])))) # (din_a[87] & (!din_b[87] $ (((!din_a[86]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_394  ) + ( Xd_0__inst_mult_7_393  ))
// Xd_0__inst_mult_7_402  = SHARE((din_a[87] & (din_b[87] & (din_a[86] & din_b[88]))))

	.dataa(!din_a[87]),
	.datab(!din_b[87]),
	.datac(!din_a[86]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_393 ),
	.sharein(Xd_0__inst_mult_7_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_400 ),
	.cout(Xd_0__inst_mult_7_401 ),
	.shareout(Xd_0__inst_mult_7_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_134 (
// Equation(s):
// Xd_0__inst_mult_4_436  = SUM(( (din_a[53] & din_b[49]) ) + ( Xd_0__inst_mult_4_430  ) + ( Xd_0__inst_mult_4_429  ))
// Xd_0__inst_mult_4_437  = CARRY(( (din_a[53] & din_b[49]) ) + ( Xd_0__inst_mult_4_430  ) + ( Xd_0__inst_mult_4_429  ))
// Xd_0__inst_mult_4_438  = SHARE((din_b[49] & din_a[54]))

	.dataa(!din_a[53]),
	.datab(!din_b[49]),
	.datac(!din_a[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_429 ),
	.sharein(Xd_0__inst_mult_4_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_436 ),
	.cout(Xd_0__inst_mult_4_437 ),
	.shareout(Xd_0__inst_mult_4_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_135 (
// Equation(s):
// Xd_0__inst_mult_4_440  = SUM(( (!din_a[51] & (((din_a[50] & din_b[52])))) # (din_a[51] & (!din_b[51] $ (((!din_a[50]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_434  ) + ( Xd_0__inst_mult_4_433  ))
// Xd_0__inst_mult_4_441  = CARRY(( (!din_a[51] & (((din_a[50] & din_b[52])))) # (din_a[51] & (!din_b[51] $ (((!din_a[50]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_434  ) + ( Xd_0__inst_mult_4_433  ))
// Xd_0__inst_mult_4_442  = SHARE((din_a[51] & (din_b[51] & (din_a[50] & din_b[52]))))

	.dataa(!din_a[51]),
	.datab(!din_b[51]),
	.datac(!din_a[50]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_433 ),
	.sharein(Xd_0__inst_mult_4_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_440 ),
	.cout(Xd_0__inst_mult_4_441 ),
	.shareout(Xd_0__inst_mult_4_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_121 (
// Equation(s):
// Xd_0__inst_mult_5_396  = SUM(( (din_a[65] & din_b[61]) ) + ( Xd_0__inst_mult_5_390  ) + ( Xd_0__inst_mult_5_389  ))
// Xd_0__inst_mult_5_397  = CARRY(( (din_a[65] & din_b[61]) ) + ( Xd_0__inst_mult_5_390  ) + ( Xd_0__inst_mult_5_389  ))
// Xd_0__inst_mult_5_398  = SHARE((din_b[61] & din_a[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[61]),
	.datac(!din_a[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_389 ),
	.sharein(Xd_0__inst_mult_5_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_396 ),
	.cout(Xd_0__inst_mult_5_397 ),
	.shareout(Xd_0__inst_mult_5_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_122 (
// Equation(s):
// Xd_0__inst_mult_5_400  = SUM(( (!din_a[63] & (((din_a[62] & din_b[64])))) # (din_a[63] & (!din_b[63] $ (((!din_a[62]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_394  ) + ( Xd_0__inst_mult_5_393  ))
// Xd_0__inst_mult_5_401  = CARRY(( (!din_a[63] & (((din_a[62] & din_b[64])))) # (din_a[63] & (!din_b[63] $ (((!din_a[62]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_394  ) + ( Xd_0__inst_mult_5_393  ))
// Xd_0__inst_mult_5_402  = SHARE((din_a[63] & (din_b[63] & (din_a[62] & din_b[64]))))

	.dataa(!din_a[63]),
	.datab(!din_b[63]),
	.datac(!din_a[62]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_393 ),
	.sharein(Xd_0__inst_mult_5_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_400 ),
	.cout(Xd_0__inst_mult_5_401 ),
	.shareout(Xd_0__inst_mult_5_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_125 (
// Equation(s):
// Xd_0__inst_mult_2_400  = SUM(( (din_a[29] & din_b[25]) ) + ( Xd_0__inst_mult_2_394  ) + ( Xd_0__inst_mult_2_393  ))
// Xd_0__inst_mult_2_401  = CARRY(( (din_a[29] & din_b[25]) ) + ( Xd_0__inst_mult_2_394  ) + ( Xd_0__inst_mult_2_393  ))
// Xd_0__inst_mult_2_402  = SHARE((din_b[25] & din_a[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[25]),
	.datac(!din_a[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_393 ),
	.sharein(Xd_0__inst_mult_2_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_400 ),
	.cout(Xd_0__inst_mult_2_401 ),
	.shareout(Xd_0__inst_mult_2_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_126 (
// Equation(s):
// Xd_0__inst_mult_2_404  = SUM(( (!din_a[27] & (((din_a[26] & din_b[28])))) # (din_a[27] & (!din_b[27] $ (((!din_a[26]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_398  ) + ( Xd_0__inst_mult_2_397  ))
// Xd_0__inst_mult_2_405  = CARRY(( (!din_a[27] & (((din_a[26] & din_b[28])))) # (din_a[27] & (!din_b[27] $ (((!din_a[26]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_398  ) + ( Xd_0__inst_mult_2_397  ))
// Xd_0__inst_mult_2_406  = SHARE((din_a[27] & (din_b[27] & (din_a[26] & din_b[28]))))

	.dataa(!din_a[27]),
	.datab(!din_b[27]),
	.datac(!din_a[26]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_397 ),
	.sharein(Xd_0__inst_mult_2_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_404 ),
	.cout(Xd_0__inst_mult_2_405 ),
	.shareout(Xd_0__inst_mult_2_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_121 (
// Equation(s):
// Xd_0__inst_mult_3_396  = SUM(( (din_a[41] & din_b[37]) ) + ( Xd_0__inst_mult_3_390  ) + ( Xd_0__inst_mult_3_389  ))
// Xd_0__inst_mult_3_397  = CARRY(( (din_a[41] & din_b[37]) ) + ( Xd_0__inst_mult_3_390  ) + ( Xd_0__inst_mult_3_389  ))
// Xd_0__inst_mult_3_398  = SHARE((din_b[37] & din_a[42]))

	.dataa(!din_a[41]),
	.datab(!din_b[37]),
	.datac(!din_a[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_389 ),
	.sharein(Xd_0__inst_mult_3_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_396 ),
	.cout(Xd_0__inst_mult_3_397 ),
	.shareout(Xd_0__inst_mult_3_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_122 (
// Equation(s):
// Xd_0__inst_mult_3_400  = SUM(( (!din_a[39] & (((din_a[38] & din_b[40])))) # (din_a[39] & (!din_b[39] $ (((!din_a[38]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_394  ) + ( Xd_0__inst_mult_3_393  ))
// Xd_0__inst_mult_3_401  = CARRY(( (!din_a[39] & (((din_a[38] & din_b[40])))) # (din_a[39] & (!din_b[39] $ (((!din_a[38]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_394  ) + ( Xd_0__inst_mult_3_393  ))
// Xd_0__inst_mult_3_402  = SHARE((din_a[39] & (din_b[39] & (din_a[38] & din_b[40]))))

	.dataa(!din_a[39]),
	.datab(!din_b[39]),
	.datac(!din_a[38]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_393 ),
	.sharein(Xd_0__inst_mult_3_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_400 ),
	.cout(Xd_0__inst_mult_3_401 ),
	.shareout(Xd_0__inst_mult_3_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_125 (
// Equation(s):
// Xd_0__inst_mult_0_400  = SUM(( (din_a[5] & din_b[1]) ) + ( Xd_0__inst_mult_0_394  ) + ( Xd_0__inst_mult_0_393  ))
// Xd_0__inst_mult_0_401  = CARRY(( (din_a[5] & din_b[1]) ) + ( Xd_0__inst_mult_0_394  ) + ( Xd_0__inst_mult_0_393  ))
// Xd_0__inst_mult_0_402  = SHARE((din_b[1] & din_a[6]))

	.dataa(!din_a[5]),
	.datab(!din_b[1]),
	.datac(!din_a[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_393 ),
	.sharein(Xd_0__inst_mult_0_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_400 ),
	.cout(Xd_0__inst_mult_0_401 ),
	.shareout(Xd_0__inst_mult_0_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_126 (
// Equation(s):
// Xd_0__inst_mult_0_404  = SUM(( (!din_a[3] & (((din_a[2] & din_b[4])))) # (din_a[3] & (!din_b[3] $ (((!din_a[2]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_398  ) + ( Xd_0__inst_mult_0_397  ))
// Xd_0__inst_mult_0_405  = CARRY(( (!din_a[3] & (((din_a[2] & din_b[4])))) # (din_a[3] & (!din_b[3] $ (((!din_a[2]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_398  ) + ( Xd_0__inst_mult_0_397  ))
// Xd_0__inst_mult_0_406  = SHARE((din_a[3] & (din_b[3] & (din_a[2] & din_b[4]))))

	.dataa(!din_a[3]),
	.datab(!din_b[3]),
	.datac(!din_a[2]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_397 ),
	.sharein(Xd_0__inst_mult_0_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_404 ),
	.cout(Xd_0__inst_mult_0_405 ),
	.shareout(Xd_0__inst_mult_0_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_125 (
// Equation(s):
// Xd_0__inst_mult_1_400  = SUM(( (din_a[17] & din_b[13]) ) + ( Xd_0__inst_mult_1_394  ) + ( Xd_0__inst_mult_1_393  ))
// Xd_0__inst_mult_1_401  = CARRY(( (din_a[17] & din_b[13]) ) + ( Xd_0__inst_mult_1_394  ) + ( Xd_0__inst_mult_1_393  ))
// Xd_0__inst_mult_1_402  = SHARE((din_b[13] & din_a[18]))

	.dataa(!din_a[17]),
	.datab(!din_b[13]),
	.datac(!din_a[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_393 ),
	.sharein(Xd_0__inst_mult_1_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_400 ),
	.cout(Xd_0__inst_mult_1_401 ),
	.shareout(Xd_0__inst_mult_1_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_126 (
// Equation(s):
// Xd_0__inst_mult_1_404  = SUM(( (!din_a[15] & (((din_a[14] & din_b[16])))) # (din_a[15] & (!din_b[15] $ (((!din_a[14]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_398  ) + ( Xd_0__inst_mult_1_397  ))
// Xd_0__inst_mult_1_405  = CARRY(( (!din_a[15] & (((din_a[14] & din_b[16])))) # (din_a[15] & (!din_b[15] $ (((!din_a[14]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_398  ) + ( Xd_0__inst_mult_1_397  ))
// Xd_0__inst_mult_1_406  = SHARE((din_a[15] & (din_b[15] & (din_a[14] & din_b[16]))))

	.dataa(!din_a[15]),
	.datab(!din_b[15]),
	.datac(!din_a[14]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_397 ),
	.sharein(Xd_0__inst_mult_1_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_404 ),
	.cout(Xd_0__inst_mult_1_405 ),
	.shareout(Xd_0__inst_mult_1_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_134 (
// Equation(s):
// Xd_0__inst_mult_12_448  = SUM(( (din_a[149] & din_b[146]) ) + ( Xd_0__inst_mult_12_442  ) + ( Xd_0__inst_mult_12_441  ))
// Xd_0__inst_mult_12_449  = CARRY(( (din_a[149] & din_b[146]) ) + ( Xd_0__inst_mult_12_442  ) + ( Xd_0__inst_mult_12_441  ))
// Xd_0__inst_mult_12_450  = SHARE((din_a[151] & din_b[145]))

	.dataa(!din_a[149]),
	.datab(!din_b[146]),
	.datac(!din_a[151]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_441 ),
	.sharein(Xd_0__inst_mult_12_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_448 ),
	.cout(Xd_0__inst_mult_12_449 ),
	.shareout(Xd_0__inst_mult_12_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_135 (
// Equation(s):
// Xd_0__inst_mult_12_452  = SUM(( (!din_a[148] & (((din_a[147] & din_b[148])))) # (din_a[148] & (!din_b[147] $ (((!din_a[147]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_446  ) + ( Xd_0__inst_mult_12_445  ))
// Xd_0__inst_mult_12_453  = CARRY(( (!din_a[148] & (((din_a[147] & din_b[148])))) # (din_a[148] & (!din_b[147] $ (((!din_a[147]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_446  ) + ( Xd_0__inst_mult_12_445  ))
// Xd_0__inst_mult_12_454  = SHARE((din_a[148] & (din_b[147] & (din_a[147] & din_b[148]))))

	.dataa(!din_a[148]),
	.datab(!din_b[147]),
	.datac(!din_a[147]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_445 ),
	.sharein(Xd_0__inst_mult_12_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_452 ),
	.cout(Xd_0__inst_mult_12_453 ),
	.shareout(Xd_0__inst_mult_12_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_131 (
// Equation(s):
// Xd_0__inst_mult_13_424  = SUM(( (din_a[161] & din_b[158]) ) + ( Xd_0__inst_mult_13_418  ) + ( Xd_0__inst_mult_13_417  ))
// Xd_0__inst_mult_13_425  = CARRY(( (din_a[161] & din_b[158]) ) + ( Xd_0__inst_mult_13_418  ) + ( Xd_0__inst_mult_13_417  ))
// Xd_0__inst_mult_13_426  = SHARE((din_a[163] & din_b[157]))

	.dataa(!din_a[161]),
	.datab(!din_b[158]),
	.datac(!din_a[163]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_417 ),
	.sharein(Xd_0__inst_mult_13_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_424 ),
	.cout(Xd_0__inst_mult_13_425 ),
	.shareout(Xd_0__inst_mult_13_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_132 (
// Equation(s):
// Xd_0__inst_mult_13_428  = SUM(( (!din_a[160] & (((din_a[159] & din_b[160])))) # (din_a[160] & (!din_b[159] $ (((!din_a[159]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_422  ) + ( Xd_0__inst_mult_13_421  ))
// Xd_0__inst_mult_13_429  = CARRY(( (!din_a[160] & (((din_a[159] & din_b[160])))) # (din_a[160] & (!din_b[159] $ (((!din_a[159]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_422  ) + ( Xd_0__inst_mult_13_421  ))
// Xd_0__inst_mult_13_430  = SHARE((din_a[160] & (din_b[159] & (din_a[159] & din_b[160]))))

	.dataa(!din_a[160]),
	.datab(!din_b[159]),
	.datac(!din_a[159]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_421 ),
	.sharein(Xd_0__inst_mult_13_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_428 ),
	.cout(Xd_0__inst_mult_13_429 ),
	.shareout(Xd_0__inst_mult_13_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_63 (
// Equation(s):
// Xd_0__inst_mult_13_63_sumout  = SUM(( (din_a[163] & din_b[156]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_64  = CARRY(( (din_a[163] & din_b[156]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_65  = SHARE(GND)

	.dataa(!din_a[163]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_13_63_sumout ),
	.cout(Xd_0__inst_mult_13_64 ),
	.shareout(Xd_0__inst_mult_13_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_135 (
// Equation(s):
// Xd_0__inst_mult_14_440  = SUM(( (din_a[173] & din_b[170]) ) + ( Xd_0__inst_mult_14_434  ) + ( Xd_0__inst_mult_14_433  ))
// Xd_0__inst_mult_14_441  = CARRY(( (din_a[173] & din_b[170]) ) + ( Xd_0__inst_mult_14_434  ) + ( Xd_0__inst_mult_14_433  ))
// Xd_0__inst_mult_14_442  = SHARE((din_a[175] & din_b[169]))

	.dataa(!din_a[173]),
	.datab(!din_b[170]),
	.datac(!din_a[175]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_433 ),
	.sharein(Xd_0__inst_mult_14_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_440 ),
	.cout(Xd_0__inst_mult_14_441 ),
	.shareout(Xd_0__inst_mult_14_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_136 (
// Equation(s):
// Xd_0__inst_mult_14_444  = SUM(( (!din_a[172] & (((din_a[171] & din_b[172])))) # (din_a[172] & (!din_b[171] $ (((!din_a[171]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_438  ) + ( Xd_0__inst_mult_14_437  ))
// Xd_0__inst_mult_14_445  = CARRY(( (!din_a[172] & (((din_a[171] & din_b[172])))) # (din_a[172] & (!din_b[171] $ (((!din_a[171]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_438  ) + ( Xd_0__inst_mult_14_437  ))
// Xd_0__inst_mult_14_446  = SHARE((din_a[172] & (din_b[171] & (din_a[171] & din_b[172]))))

	.dataa(!din_a[172]),
	.datab(!din_b[171]),
	.datac(!din_a[171]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_437 ),
	.sharein(Xd_0__inst_mult_14_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_444 ),
	.cout(Xd_0__inst_mult_14_445 ),
	.shareout(Xd_0__inst_mult_14_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_138 (
// Equation(s):
// Xd_0__inst_mult_15_452  = SUM(( (din_a[185] & din_b[182]) ) + ( Xd_0__inst_mult_15_446  ) + ( Xd_0__inst_mult_15_445  ))
// Xd_0__inst_mult_15_453  = CARRY(( (din_a[185] & din_b[182]) ) + ( Xd_0__inst_mult_15_446  ) + ( Xd_0__inst_mult_15_445  ))
// Xd_0__inst_mult_15_454  = SHARE((din_a[187] & din_b[181]))

	.dataa(!din_a[185]),
	.datab(!din_b[182]),
	.datac(!din_a[187]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_445 ),
	.sharein(Xd_0__inst_mult_15_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_452 ),
	.cout(Xd_0__inst_mult_15_453 ),
	.shareout(Xd_0__inst_mult_15_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_139 (
// Equation(s):
// Xd_0__inst_mult_15_456  = SUM(( (!din_a[184] & (((din_a[183] & din_b[184])))) # (din_a[184] & (!din_b[183] $ (((!din_a[183]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_450  ) + ( Xd_0__inst_mult_15_449  ))
// Xd_0__inst_mult_15_457  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[184])))) # (din_a[184] & (!din_b[183] $ (((!din_a[183]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_450  ) + ( Xd_0__inst_mult_15_449  ))
// Xd_0__inst_mult_15_458  = SHARE((din_a[184] & (din_b[183] & (din_a[183] & din_b[184]))))

	.dataa(!din_a[184]),
	.datab(!din_b[183]),
	.datac(!din_a[183]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_449 ),
	.sharein(Xd_0__inst_mult_15_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_456 ),
	.cout(Xd_0__inst_mult_15_457 ),
	.shareout(Xd_0__inst_mult_15_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_127 (
// Equation(s):
// Xd_0__inst_mult_10_420  = SUM(( (din_a[125] & din_b[122]) ) + ( Xd_0__inst_mult_10_414  ) + ( Xd_0__inst_mult_10_413  ))
// Xd_0__inst_mult_10_421  = CARRY(( (din_a[125] & din_b[122]) ) + ( Xd_0__inst_mult_10_414  ) + ( Xd_0__inst_mult_10_413  ))
// Xd_0__inst_mult_10_422  = SHARE((din_a[127] & din_b[121]))

	.dataa(!din_a[125]),
	.datab(!din_b[122]),
	.datac(!din_a[127]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_413 ),
	.sharein(Xd_0__inst_mult_10_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_420 ),
	.cout(Xd_0__inst_mult_10_421 ),
	.shareout(Xd_0__inst_mult_10_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_128 (
// Equation(s):
// Xd_0__inst_mult_10_424  = SUM(( (!din_a[124] & (((din_a[123] & din_b[124])))) # (din_a[124] & (!din_b[123] $ (((!din_a[123]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_418  ) + ( Xd_0__inst_mult_10_417  ))
// Xd_0__inst_mult_10_425  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[124])))) # (din_a[124] & (!din_b[123] $ (((!din_a[123]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_418  ) + ( Xd_0__inst_mult_10_417  ))
// Xd_0__inst_mult_10_426  = SHARE((din_a[124] & (din_b[123] & (din_a[123] & din_b[124]))))

	.dataa(!din_a[124]),
	.datab(!din_b[123]),
	.datac(!din_a[123]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_417 ),
	.sharein(Xd_0__inst_mult_10_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_424 ),
	.cout(Xd_0__inst_mult_10_425 ),
	.shareout(Xd_0__inst_mult_10_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_131 (
// Equation(s):
// Xd_0__inst_mult_11_424  = SUM(( (din_a[137] & din_b[134]) ) + ( Xd_0__inst_mult_11_418  ) + ( Xd_0__inst_mult_11_417  ))
// Xd_0__inst_mult_11_425  = CARRY(( (din_a[137] & din_b[134]) ) + ( Xd_0__inst_mult_11_418  ) + ( Xd_0__inst_mult_11_417  ))
// Xd_0__inst_mult_11_426  = SHARE((din_a[139] & din_b[133]))

	.dataa(!din_a[137]),
	.datab(!din_b[134]),
	.datac(!din_a[139]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_417 ),
	.sharein(Xd_0__inst_mult_11_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_424 ),
	.cout(Xd_0__inst_mult_11_425 ),
	.shareout(Xd_0__inst_mult_11_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_132 (
// Equation(s):
// Xd_0__inst_mult_11_428  = SUM(( (!din_a[136] & (((din_a[135] & din_b[136])))) # (din_a[136] & (!din_b[135] $ (((!din_a[135]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_422  ) + ( Xd_0__inst_mult_11_421  ))
// Xd_0__inst_mult_11_429  = CARRY(( (!din_a[136] & (((din_a[135] & din_b[136])))) # (din_a[136] & (!din_b[135] $ (((!din_a[135]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_422  ) + ( Xd_0__inst_mult_11_421  ))
// Xd_0__inst_mult_11_430  = SHARE((din_a[136] & (din_b[135] & (din_a[135] & din_b[136]))))

	.dataa(!din_a[136]),
	.datab(!din_b[135]),
	.datac(!din_a[135]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_421 ),
	.sharein(Xd_0__inst_mult_11_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_428 ),
	.cout(Xd_0__inst_mult_11_429 ),
	.shareout(Xd_0__inst_mult_11_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_63 (
// Equation(s):
// Xd_0__inst_mult_11_63_sumout  = SUM(( (din_a[139] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_64  = CARRY(( (din_a[139] & din_b[132]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_65  = SHARE(GND)

	.dataa(!din_a[139]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_63_sumout ),
	.cout(Xd_0__inst_mult_11_64 ),
	.shareout(Xd_0__inst_mult_11_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_131 (
// Equation(s):
// Xd_0__inst_mult_8_424  = SUM(( (din_a[101] & din_b[98]) ) + ( Xd_0__inst_mult_8_418  ) + ( Xd_0__inst_mult_8_417  ))
// Xd_0__inst_mult_8_425  = CARRY(( (din_a[101] & din_b[98]) ) + ( Xd_0__inst_mult_8_418  ) + ( Xd_0__inst_mult_8_417  ))
// Xd_0__inst_mult_8_426  = SHARE((din_a[103] & din_b[97]))

	.dataa(!din_a[101]),
	.datab(!din_b[98]),
	.datac(!din_a[103]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_417 ),
	.sharein(Xd_0__inst_mult_8_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_424 ),
	.cout(Xd_0__inst_mult_8_425 ),
	.shareout(Xd_0__inst_mult_8_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_132 (
// Equation(s):
// Xd_0__inst_mult_8_428  = SUM(( (!din_a[100] & (((din_a[99] & din_b[100])))) # (din_a[100] & (!din_b[99] $ (((!din_a[99]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_422  ) + ( Xd_0__inst_mult_8_421  ))
// Xd_0__inst_mult_8_429  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[100])))) # (din_a[100] & (!din_b[99] $ (((!din_a[99]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_422  ) + ( Xd_0__inst_mult_8_421  ))
// Xd_0__inst_mult_8_430  = SHARE((din_a[100] & (din_b[99] & (din_a[99] & din_b[100]))))

	.dataa(!din_a[100]),
	.datab(!din_b[99]),
	.datac(!din_a[99]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_421 ),
	.sharein(Xd_0__inst_mult_8_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_428 ),
	.cout(Xd_0__inst_mult_8_429 ),
	.shareout(Xd_0__inst_mult_8_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_63 (
// Equation(s):
// Xd_0__inst_mult_8_63_sumout  = SUM(( (din_a[103] & din_b[96]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_64  = CARRY(( (din_a[103] & din_b[96]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_65  = SHARE(GND)

	.dataa(!din_a[103]),
	.datab(!din_b[96]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_8_63_sumout ),
	.cout(Xd_0__inst_mult_8_64 ),
	.shareout(Xd_0__inst_mult_8_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_127 (
// Equation(s):
// Xd_0__inst_mult_9_420  = SUM(( (din_a[113] & din_b[110]) ) + ( Xd_0__inst_mult_9_414  ) + ( Xd_0__inst_mult_9_413  ))
// Xd_0__inst_mult_9_421  = CARRY(( (din_a[113] & din_b[110]) ) + ( Xd_0__inst_mult_9_414  ) + ( Xd_0__inst_mult_9_413  ))
// Xd_0__inst_mult_9_422  = SHARE((din_a[115] & din_b[109]))

	.dataa(!din_a[113]),
	.datab(!din_b[110]),
	.datac(!din_a[115]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_413 ),
	.sharein(Xd_0__inst_mult_9_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_420 ),
	.cout(Xd_0__inst_mult_9_421 ),
	.shareout(Xd_0__inst_mult_9_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_128 (
// Equation(s):
// Xd_0__inst_mult_9_424  = SUM(( (!din_a[112] & (((din_a[111] & din_b[112])))) # (din_a[112] & (!din_b[111] $ (((!din_a[111]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_418  ) + ( Xd_0__inst_mult_9_417  ))
// Xd_0__inst_mult_9_425  = CARRY(( (!din_a[112] & (((din_a[111] & din_b[112])))) # (din_a[112] & (!din_b[111] $ (((!din_a[111]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_418  ) + ( Xd_0__inst_mult_9_417  ))
// Xd_0__inst_mult_9_426  = SHARE((din_a[112] & (din_b[111] & (din_a[111] & din_b[112]))))

	.dataa(!din_a[112]),
	.datab(!din_b[111]),
	.datac(!din_a[111]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_417 ),
	.sharein(Xd_0__inst_mult_9_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_424 ),
	.cout(Xd_0__inst_mult_9_425 ),
	.shareout(Xd_0__inst_mult_9_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_59 (
// Equation(s):
// Xd_0__inst_mult_9_59_sumout  = SUM(( (din_a[115] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_60  = CARRY(( (din_a[115] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_61  = SHARE(GND)

	.dataa(!din_a[115]),
	.datab(!din_b[108]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_59_sumout ),
	.cout(Xd_0__inst_mult_9_60 ),
	.shareout(Xd_0__inst_mult_9_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_127 (
// Equation(s):
// Xd_0__inst_mult_6_420  = SUM(( (din_a[77] & din_b[74]) ) + ( Xd_0__inst_mult_6_414  ) + ( Xd_0__inst_mult_6_413  ))
// Xd_0__inst_mult_6_421  = CARRY(( (din_a[77] & din_b[74]) ) + ( Xd_0__inst_mult_6_414  ) + ( Xd_0__inst_mult_6_413  ))
// Xd_0__inst_mult_6_422  = SHARE((din_a[79] & din_b[73]))

	.dataa(!din_a[77]),
	.datab(!din_b[74]),
	.datac(!din_a[79]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_413 ),
	.sharein(Xd_0__inst_mult_6_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_420 ),
	.cout(Xd_0__inst_mult_6_421 ),
	.shareout(Xd_0__inst_mult_6_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_128 (
// Equation(s):
// Xd_0__inst_mult_6_424  = SUM(( (!din_a[76] & (((din_a[75] & din_b[76])))) # (din_a[76] & (!din_b[75] $ (((!din_a[75]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_418  ) + ( Xd_0__inst_mult_6_417  ))
// Xd_0__inst_mult_6_425  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[76])))) # (din_a[76] & (!din_b[75] $ (((!din_a[75]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_418  ) + ( Xd_0__inst_mult_6_417  ))
// Xd_0__inst_mult_6_426  = SHARE((din_a[76] & (din_b[75] & (din_a[75] & din_b[76]))))

	.dataa(!din_a[76]),
	.datab(!din_b[75]),
	.datac(!din_a[75]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_417 ),
	.sharein(Xd_0__inst_mult_6_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_424 ),
	.cout(Xd_0__inst_mult_6_425 ),
	.shareout(Xd_0__inst_mult_6_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_59 (
// Equation(s):
// Xd_0__inst_mult_6_59_sumout  = SUM(( (din_a[79] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_60  = CARRY(( (din_a[79] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_61  = SHARE(GND)

	.dataa(!din_a[79]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_59_sumout ),
	.cout(Xd_0__inst_mult_6_60 ),
	.shareout(Xd_0__inst_mult_6_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_123 (
// Equation(s):
// Xd_0__inst_mult_7_404  = SUM(( (din_a[89] & din_b[86]) ) + ( Xd_0__inst_mult_7_398  ) + ( Xd_0__inst_mult_7_397  ))
// Xd_0__inst_mult_7_405  = CARRY(( (din_a[89] & din_b[86]) ) + ( Xd_0__inst_mult_7_398  ) + ( Xd_0__inst_mult_7_397  ))
// Xd_0__inst_mult_7_406  = SHARE((din_a[91] & din_b[85]))

	.dataa(!din_a[89]),
	.datab(!din_b[86]),
	.datac(!din_a[91]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_397 ),
	.sharein(Xd_0__inst_mult_7_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_404 ),
	.cout(Xd_0__inst_mult_7_405 ),
	.shareout(Xd_0__inst_mult_7_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_124 (
// Equation(s):
// Xd_0__inst_mult_7_408  = SUM(( (!din_a[88] & (((din_a[87] & din_b[88])))) # (din_a[88] & (!din_b[87] $ (((!din_a[87]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_402  ) + ( Xd_0__inst_mult_7_401  ))
// Xd_0__inst_mult_7_409  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[88])))) # (din_a[88] & (!din_b[87] $ (((!din_a[87]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_402  ) + ( Xd_0__inst_mult_7_401  ))
// Xd_0__inst_mult_7_410  = SHARE((din_a[88] & (din_b[87] & (din_a[87] & din_b[88]))))

	.dataa(!din_a[88]),
	.datab(!din_b[87]),
	.datac(!din_a[87]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_401 ),
	.sharein(Xd_0__inst_mult_7_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_408 ),
	.cout(Xd_0__inst_mult_7_409 ),
	.shareout(Xd_0__inst_mult_7_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_55 (
// Equation(s):
// Xd_0__inst_mult_7_55_sumout  = SUM(( (din_a[91] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_56  = CARRY(( (din_a[91] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_57  = SHARE(GND)

	.dataa(!din_a[91]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_55_sumout ),
	.cout(Xd_0__inst_mult_7_56 ),
	.shareout(Xd_0__inst_mult_7_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_136 (
// Equation(s):
// Xd_0__inst_mult_4_444  = SUM(( (din_a[53] & din_b[50]) ) + ( Xd_0__inst_mult_4_438  ) + ( Xd_0__inst_mult_4_437  ))
// Xd_0__inst_mult_4_445  = CARRY(( (din_a[53] & din_b[50]) ) + ( Xd_0__inst_mult_4_438  ) + ( Xd_0__inst_mult_4_437  ))
// Xd_0__inst_mult_4_446  = SHARE((din_a[55] & din_b[49]))

	.dataa(!din_a[53]),
	.datab(!din_b[50]),
	.datac(!din_a[55]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_437 ),
	.sharein(Xd_0__inst_mult_4_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_444 ),
	.cout(Xd_0__inst_mult_4_445 ),
	.shareout(Xd_0__inst_mult_4_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_137 (
// Equation(s):
// Xd_0__inst_mult_4_448  = SUM(( (!din_a[52] & (((din_a[51] & din_b[52])))) # (din_a[52] & (!din_b[51] $ (((!din_a[51]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_442  ) + ( Xd_0__inst_mult_4_441  ))
// Xd_0__inst_mult_4_449  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[52])))) # (din_a[52] & (!din_b[51] $ (((!din_a[51]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_442  ) + ( Xd_0__inst_mult_4_441  ))
// Xd_0__inst_mult_4_450  = SHARE((din_a[52] & (din_b[51] & (din_a[51] & din_b[52]))))

	.dataa(!din_a[52]),
	.datab(!din_b[51]),
	.datac(!din_a[51]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_441 ),
	.sharein(Xd_0__inst_mult_4_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_448 ),
	.cout(Xd_0__inst_mult_4_449 ),
	.shareout(Xd_0__inst_mult_4_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_59 (
// Equation(s):
// Xd_0__inst_mult_4_59_sumout  = SUM(( (din_a[55] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_60  = CARRY(( (din_a[55] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_61  = SHARE(GND)

	.dataa(!din_a[55]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_59_sumout ),
	.cout(Xd_0__inst_mult_4_60 ),
	.shareout(Xd_0__inst_mult_4_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_123 (
// Equation(s):
// Xd_0__inst_mult_5_404  = SUM(( (din_a[65] & din_b[62]) ) + ( Xd_0__inst_mult_5_398  ) + ( Xd_0__inst_mult_5_397  ))
// Xd_0__inst_mult_5_405  = CARRY(( (din_a[65] & din_b[62]) ) + ( Xd_0__inst_mult_5_398  ) + ( Xd_0__inst_mult_5_397  ))
// Xd_0__inst_mult_5_406  = SHARE((din_a[67] & din_b[61]))

	.dataa(!din_a[65]),
	.datab(!din_b[62]),
	.datac(!din_a[67]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_397 ),
	.sharein(Xd_0__inst_mult_5_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_404 ),
	.cout(Xd_0__inst_mult_5_405 ),
	.shareout(Xd_0__inst_mult_5_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_124 (
// Equation(s):
// Xd_0__inst_mult_5_408  = SUM(( (!din_a[64] & (((din_a[63] & din_b[64])))) # (din_a[64] & (!din_b[63] $ (((!din_a[63]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_402  ) + ( Xd_0__inst_mult_5_401  ))
// Xd_0__inst_mult_5_409  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[64])))) # (din_a[64] & (!din_b[63] $ (((!din_a[63]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_402  ) + ( Xd_0__inst_mult_5_401  ))
// Xd_0__inst_mult_5_410  = SHARE((din_a[64] & (din_b[63] & (din_a[63] & din_b[64]))))

	.dataa(!din_a[64]),
	.datab(!din_b[63]),
	.datac(!din_a[63]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_401 ),
	.sharein(Xd_0__inst_mult_5_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_408 ),
	.cout(Xd_0__inst_mult_5_409 ),
	.shareout(Xd_0__inst_mult_5_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_59 (
// Equation(s):
// Xd_0__inst_mult_5_59_sumout  = SUM(( (din_a[67] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_60  = CARRY(( (din_a[67] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_61  = SHARE(GND)

	.dataa(!din_a[67]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_59_sumout ),
	.cout(Xd_0__inst_mult_5_60 ),
	.shareout(Xd_0__inst_mult_5_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_127 (
// Equation(s):
// Xd_0__inst_mult_2_408  = SUM(( (din_a[29] & din_b[26]) ) + ( Xd_0__inst_mult_2_402  ) + ( Xd_0__inst_mult_2_401  ))
// Xd_0__inst_mult_2_409  = CARRY(( (din_a[29] & din_b[26]) ) + ( Xd_0__inst_mult_2_402  ) + ( Xd_0__inst_mult_2_401  ))
// Xd_0__inst_mult_2_410  = SHARE((din_a[31] & din_b[25]))

	.dataa(!din_a[29]),
	.datab(!din_b[26]),
	.datac(!din_a[31]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_401 ),
	.sharein(Xd_0__inst_mult_2_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_408 ),
	.cout(Xd_0__inst_mult_2_409 ),
	.shareout(Xd_0__inst_mult_2_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_128 (
// Equation(s):
// Xd_0__inst_mult_2_412  = SUM(( (!din_a[28] & (((din_a[27] & din_b[28])))) # (din_a[28] & (!din_b[27] $ (((!din_a[27]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_406  ) + ( Xd_0__inst_mult_2_405  ))
// Xd_0__inst_mult_2_413  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[28])))) # (din_a[28] & (!din_b[27] $ (((!din_a[27]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_406  ) + ( Xd_0__inst_mult_2_405  ))
// Xd_0__inst_mult_2_414  = SHARE((din_a[28] & (din_b[27] & (din_a[27] & din_b[28]))))

	.dataa(!din_a[28]),
	.datab(!din_b[27]),
	.datac(!din_a[27]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_405 ),
	.sharein(Xd_0__inst_mult_2_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_412 ),
	.cout(Xd_0__inst_mult_2_413 ),
	.shareout(Xd_0__inst_mult_2_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_123 (
// Equation(s):
// Xd_0__inst_mult_3_404  = SUM(( (din_a[41] & din_b[38]) ) + ( Xd_0__inst_mult_3_398  ) + ( Xd_0__inst_mult_3_397  ))
// Xd_0__inst_mult_3_405  = CARRY(( (din_a[41] & din_b[38]) ) + ( Xd_0__inst_mult_3_398  ) + ( Xd_0__inst_mult_3_397  ))
// Xd_0__inst_mult_3_406  = SHARE((din_a[43] & din_b[37]))

	.dataa(!din_a[41]),
	.datab(!din_b[38]),
	.datac(!din_a[43]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_397 ),
	.sharein(Xd_0__inst_mult_3_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_404 ),
	.cout(Xd_0__inst_mult_3_405 ),
	.shareout(Xd_0__inst_mult_3_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_124 (
// Equation(s):
// Xd_0__inst_mult_3_408  = SUM(( (!din_a[40] & (((din_a[39] & din_b[40])))) # (din_a[40] & (!din_b[39] $ (((!din_a[39]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_402  ) + ( Xd_0__inst_mult_3_401  ))
// Xd_0__inst_mult_3_409  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[40])))) # (din_a[40] & (!din_b[39] $ (((!din_a[39]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_402  ) + ( Xd_0__inst_mult_3_401  ))
// Xd_0__inst_mult_3_410  = SHARE((din_a[40] & (din_b[39] & (din_a[39] & din_b[40]))))

	.dataa(!din_a[40]),
	.datab(!din_b[39]),
	.datac(!din_a[39]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_401 ),
	.sharein(Xd_0__inst_mult_3_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_408 ),
	.cout(Xd_0__inst_mult_3_409 ),
	.shareout(Xd_0__inst_mult_3_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_127 (
// Equation(s):
// Xd_0__inst_mult_0_408  = SUM(( (din_a[5] & din_b[2]) ) + ( Xd_0__inst_mult_0_402  ) + ( Xd_0__inst_mult_0_401  ))
// Xd_0__inst_mult_0_409  = CARRY(( (din_a[5] & din_b[2]) ) + ( Xd_0__inst_mult_0_402  ) + ( Xd_0__inst_mult_0_401  ))
// Xd_0__inst_mult_0_410  = SHARE((din_a[7] & din_b[1]))

	.dataa(!din_a[5]),
	.datab(!din_b[2]),
	.datac(!din_a[7]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_401 ),
	.sharein(Xd_0__inst_mult_0_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_408 ),
	.cout(Xd_0__inst_mult_0_409 ),
	.shareout(Xd_0__inst_mult_0_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_128 (
// Equation(s):
// Xd_0__inst_mult_0_412  = SUM(( (!din_a[4] & (((din_a[3] & din_b[4])))) # (din_a[4] & (!din_b[3] $ (((!din_a[3]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_406  ) + ( Xd_0__inst_mult_0_405  ))
// Xd_0__inst_mult_0_413  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[4])))) # (din_a[4] & (!din_b[3] $ (((!din_a[3]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_406  ) + ( Xd_0__inst_mult_0_405  ))
// Xd_0__inst_mult_0_414  = SHARE((din_a[4] & (din_b[3] & (din_a[3] & din_b[4]))))

	.dataa(!din_a[4]),
	.datab(!din_b[3]),
	.datac(!din_a[3]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_405 ),
	.sharein(Xd_0__inst_mult_0_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_412 ),
	.cout(Xd_0__inst_mult_0_413 ),
	.shareout(Xd_0__inst_mult_0_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_127 (
// Equation(s):
// Xd_0__inst_mult_1_408  = SUM(( (din_a[17] & din_b[14]) ) + ( Xd_0__inst_mult_1_402  ) + ( Xd_0__inst_mult_1_401  ))
// Xd_0__inst_mult_1_409  = CARRY(( (din_a[17] & din_b[14]) ) + ( Xd_0__inst_mult_1_402  ) + ( Xd_0__inst_mult_1_401  ))
// Xd_0__inst_mult_1_410  = SHARE((din_a[19] & din_b[13]))

	.dataa(!din_a[17]),
	.datab(!din_b[14]),
	.datac(!din_a[19]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_401 ),
	.sharein(Xd_0__inst_mult_1_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_408 ),
	.cout(Xd_0__inst_mult_1_409 ),
	.shareout(Xd_0__inst_mult_1_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_128 (
// Equation(s):
// Xd_0__inst_mult_1_412  = SUM(( (!din_a[16] & (((din_a[15] & din_b[16])))) # (din_a[16] & (!din_b[15] $ (((!din_a[15]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_406  ) + ( Xd_0__inst_mult_1_405  ))
// Xd_0__inst_mult_1_413  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[16])))) # (din_a[16] & (!din_b[15] $ (((!din_a[15]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_406  ) + ( Xd_0__inst_mult_1_405  ))
// Xd_0__inst_mult_1_414  = SHARE((din_a[16] & (din_b[15] & (din_a[15] & din_b[16]))))

	.dataa(!din_a[16]),
	.datab(!din_b[15]),
	.datac(!din_a[15]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_405 ),
	.sharein(Xd_0__inst_mult_1_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_412 ),
	.cout(Xd_0__inst_mult_1_413 ),
	.shareout(Xd_0__inst_mult_1_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_136 (
// Equation(s):
// Xd_0__inst_mult_12_456  = SUM(( (din_a[150] & din_b[146]) ) + ( Xd_0__inst_mult_12_450  ) + ( Xd_0__inst_mult_12_449  ))
// Xd_0__inst_mult_12_457  = CARRY(( (din_a[150] & din_b[146]) ) + ( Xd_0__inst_mult_12_450  ) + ( Xd_0__inst_mult_12_449  ))
// Xd_0__inst_mult_12_458  = SHARE((din_a[152] & din_b[145]))

	.dataa(!din_a[150]),
	.datab(!din_b[146]),
	.datac(!din_a[152]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_449 ),
	.sharein(Xd_0__inst_mult_12_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_456 ),
	.cout(Xd_0__inst_mult_12_457 ),
	.shareout(Xd_0__inst_mult_12_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_137 (
// Equation(s):
// Xd_0__inst_mult_12_460  = SUM(( (!din_a[149] & (((din_a[148] & din_b[148])))) # (din_a[149] & (!din_b[147] $ (((!din_a[148]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_454  ) + ( Xd_0__inst_mult_12_453  ))
// Xd_0__inst_mult_12_461  = CARRY(( (!din_a[149] & (((din_a[148] & din_b[148])))) # (din_a[149] & (!din_b[147] $ (((!din_a[148]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_454  ) + ( Xd_0__inst_mult_12_453  ))
// Xd_0__inst_mult_12_462  = SHARE((din_a[149] & (din_b[147] & (din_a[148] & din_b[148]))))

	.dataa(!din_a[149]),
	.datab(!din_b[147]),
	.datac(!din_a[148]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_453 ),
	.sharein(Xd_0__inst_mult_12_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_460 ),
	.cout(Xd_0__inst_mult_12_461 ),
	.shareout(Xd_0__inst_mult_12_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_138 (
// Equation(s):
// Xd_0__inst_mult_12_464  = SUM(( (!din_a[146] & (((din_a[147] & din_b[149])))) # (din_a[146] & (!din_b[150] $ (((!din_a[147]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_12_338  ) + ( Xd_0__inst_mult_12_337  ))
// Xd_0__inst_mult_12_465  = CARRY(( (!din_a[146] & (((din_a[147] & din_b[149])))) # (din_a[146] & (!din_b[150] $ (((!din_a[147]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_12_338  ) + ( Xd_0__inst_mult_12_337  ))
// Xd_0__inst_mult_12_466  = SHARE((din_a[146] & (din_b[150] & (din_a[147] & din_b[149]))))

	.dataa(!din_a[146]),
	.datab(!din_b[150]),
	.datac(!din_a[147]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_337 ),
	.sharein(Xd_0__inst_mult_12_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_464 ),
	.cout(Xd_0__inst_mult_12_465 ),
	.shareout(Xd_0__inst_mult_12_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_139 (
// Equation(s):
// Xd_0__inst_mult_12_469  = CARRY(( GND ) + ( Xd_0__inst_i29_31  ) + ( Xd_0__inst_i29_30  ))
// Xd_0__inst_mult_12_470  = SHARE((din_a[144] & din_b[152]))

	.dataa(!din_a[144]),
	.datab(!din_b[152]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_30 ),
	.sharein(Xd_0__inst_i29_31 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_469 ),
	.shareout(Xd_0__inst_mult_12_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_133 (
// Equation(s):
// Xd_0__inst_mult_13_432  = SUM(( (din_a[162] & din_b[158]) ) + ( Xd_0__inst_mult_13_426  ) + ( Xd_0__inst_mult_13_425  ))
// Xd_0__inst_mult_13_433  = CARRY(( (din_a[162] & din_b[158]) ) + ( Xd_0__inst_mult_13_426  ) + ( Xd_0__inst_mult_13_425  ))
// Xd_0__inst_mult_13_434  = SHARE((din_a[164] & din_b[157]))

	.dataa(!din_a[162]),
	.datab(!din_b[158]),
	.datac(!din_a[164]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_425 ),
	.sharein(Xd_0__inst_mult_13_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_432 ),
	.cout(Xd_0__inst_mult_13_433 ),
	.shareout(Xd_0__inst_mult_13_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_134 (
// Equation(s):
// Xd_0__inst_mult_13_436  = SUM(( (!din_a[161] & (((din_a[160] & din_b[160])))) # (din_a[161] & (!din_b[159] $ (((!din_a[160]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_430  ) + ( Xd_0__inst_mult_13_429  ))
// Xd_0__inst_mult_13_437  = CARRY(( (!din_a[161] & (((din_a[160] & din_b[160])))) # (din_a[161] & (!din_b[159] $ (((!din_a[160]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_430  ) + ( Xd_0__inst_mult_13_429  ))
// Xd_0__inst_mult_13_438  = SHARE((din_a[161] & (din_b[159] & (din_a[160] & din_b[160]))))

	.dataa(!din_a[161]),
	.datab(!din_b[159]),
	.datac(!din_a[160]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_429 ),
	.sharein(Xd_0__inst_mult_13_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_436 ),
	.cout(Xd_0__inst_mult_13_437 ),
	.shareout(Xd_0__inst_mult_13_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_135 (
// Equation(s):
// Xd_0__inst_mult_13_440  = SUM(( (!din_a[158] & (((din_a[159] & din_b[161])))) # (din_a[158] & (!din_b[162] $ (((!din_a[159]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_13_318  ) + ( Xd_0__inst_mult_13_317  ))
// Xd_0__inst_mult_13_441  = CARRY(( (!din_a[158] & (((din_a[159] & din_b[161])))) # (din_a[158] & (!din_b[162] $ (((!din_a[159]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_13_318  ) + ( Xd_0__inst_mult_13_317  ))
// Xd_0__inst_mult_13_442  = SHARE((din_a[158] & (din_b[162] & (din_a[159] & din_b[161]))))

	.dataa(!din_a[158]),
	.datab(!din_b[162]),
	.datac(!din_a[159]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_317 ),
	.sharein(Xd_0__inst_mult_13_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_440 ),
	.cout(Xd_0__inst_mult_13_441 ),
	.shareout(Xd_0__inst_mult_13_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_136 (
// Equation(s):
// Xd_0__inst_mult_13_445  = CARRY(( GND ) + ( Xd_0__inst_i29_15  ) + ( Xd_0__inst_i29_14  ))
// Xd_0__inst_mult_13_446  = SHARE((din_a[156] & din_b[164]))

	.dataa(!din_a[156]),
	.datab(!din_b[164]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_14 ),
	.sharein(Xd_0__inst_i29_15 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_445 ),
	.shareout(Xd_0__inst_mult_13_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_137 (
// Equation(s):
// Xd_0__inst_mult_14_448  = SUM(( (din_a[174] & din_b[170]) ) + ( Xd_0__inst_mult_14_442  ) + ( Xd_0__inst_mult_14_441  ))
// Xd_0__inst_mult_14_449  = CARRY(( (din_a[174] & din_b[170]) ) + ( Xd_0__inst_mult_14_442  ) + ( Xd_0__inst_mult_14_441  ))
// Xd_0__inst_mult_14_450  = SHARE((din_a[176] & din_b[169]))

	.dataa(!din_a[174]),
	.datab(!din_b[170]),
	.datac(!din_a[176]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_441 ),
	.sharein(Xd_0__inst_mult_14_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_448 ),
	.cout(Xd_0__inst_mult_14_449 ),
	.shareout(Xd_0__inst_mult_14_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_138 (
// Equation(s):
// Xd_0__inst_mult_14_452  = SUM(( (!din_a[173] & (((din_a[172] & din_b[172])))) # (din_a[173] & (!din_b[171] $ (((!din_a[172]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_446  ) + ( Xd_0__inst_mult_14_445  ))
// Xd_0__inst_mult_14_453  = CARRY(( (!din_a[173] & (((din_a[172] & din_b[172])))) # (din_a[173] & (!din_b[171] $ (((!din_a[172]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_446  ) + ( Xd_0__inst_mult_14_445  ))
// Xd_0__inst_mult_14_454  = SHARE((din_a[173] & (din_b[171] & (din_a[172] & din_b[172]))))

	.dataa(!din_a[173]),
	.datab(!din_b[171]),
	.datac(!din_a[172]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_445 ),
	.sharein(Xd_0__inst_mult_14_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_452 ),
	.cout(Xd_0__inst_mult_14_453 ),
	.shareout(Xd_0__inst_mult_14_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_139 (
// Equation(s):
// Xd_0__inst_mult_14_456  = SUM(( (!din_a[170] & (((din_a[171] & din_b[173])))) # (din_a[170] & (!din_b[174] $ (((!din_a[171]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_14_342  ) + ( Xd_0__inst_mult_14_341  ))
// Xd_0__inst_mult_14_457  = CARRY(( (!din_a[170] & (((din_a[171] & din_b[173])))) # (din_a[170] & (!din_b[174] $ (((!din_a[171]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_14_342  ) + ( Xd_0__inst_mult_14_341  ))
// Xd_0__inst_mult_14_458  = SHARE((din_a[170] & (din_b[174] & (din_a[171] & din_b[173]))))

	.dataa(!din_a[170]),
	.datab(!din_b[174]),
	.datac(!din_a[171]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_341 ),
	.sharein(Xd_0__inst_mult_14_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_456 ),
	.cout(Xd_0__inst_mult_14_457 ),
	.shareout(Xd_0__inst_mult_14_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_140 (
// Equation(s):
// Xd_0__inst_mult_14_461  = CARRY(( GND ) + ( Xd_0__inst_mult_10_45  ) + ( Xd_0__inst_mult_10_44  ))
// Xd_0__inst_mult_14_462  = SHARE((din_a[168] & din_b[176]))

	.dataa(!din_a[168]),
	.datab(!din_b[176]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_44 ),
	.sharein(Xd_0__inst_mult_10_45 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_461 ),
	.shareout(Xd_0__inst_mult_14_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_140 (
// Equation(s):
// Xd_0__inst_mult_15_460  = SUM(( (din_a[186] & din_b[182]) ) + ( Xd_0__inst_mult_15_454  ) + ( Xd_0__inst_mult_15_453  ))
// Xd_0__inst_mult_15_461  = CARRY(( (din_a[186] & din_b[182]) ) + ( Xd_0__inst_mult_15_454  ) + ( Xd_0__inst_mult_15_453  ))
// Xd_0__inst_mult_15_462  = SHARE((din_a[188] & din_b[181]))

	.dataa(!din_a[186]),
	.datab(!din_b[182]),
	.datac(!din_a[188]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_453 ),
	.sharein(Xd_0__inst_mult_15_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_460 ),
	.cout(Xd_0__inst_mult_15_461 ),
	.shareout(Xd_0__inst_mult_15_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_141 (
// Equation(s):
// Xd_0__inst_mult_15_464  = SUM(( (!din_a[185] & (((din_a[184] & din_b[184])))) # (din_a[185] & (!din_b[183] $ (((!din_a[184]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_458  ) + ( Xd_0__inst_mult_15_457  ))
// Xd_0__inst_mult_15_465  = CARRY(( (!din_a[185] & (((din_a[184] & din_b[184])))) # (din_a[185] & (!din_b[183] $ (((!din_a[184]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_458  ) + ( Xd_0__inst_mult_15_457  ))
// Xd_0__inst_mult_15_466  = SHARE((din_a[185] & (din_b[183] & (din_a[184] & din_b[184]))))

	.dataa(!din_a[185]),
	.datab(!din_b[183]),
	.datac(!din_a[184]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_457 ),
	.sharein(Xd_0__inst_mult_15_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_464 ),
	.cout(Xd_0__inst_mult_15_465 ),
	.shareout(Xd_0__inst_mult_15_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_142 (
// Equation(s):
// Xd_0__inst_mult_15_468  = SUM(( (!din_a[182] & (((din_a[183] & din_b[185])))) # (din_a[182] & (!din_b[186] $ (((!din_a[183]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_15_342  ) + ( Xd_0__inst_mult_15_341  ))
// Xd_0__inst_mult_15_469  = CARRY(( (!din_a[182] & (((din_a[183] & din_b[185])))) # (din_a[182] & (!din_b[186] $ (((!din_a[183]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_15_342  ) + ( Xd_0__inst_mult_15_341  ))
// Xd_0__inst_mult_15_470  = SHARE((din_a[182] & (din_b[186] & (din_a[183] & din_b[185]))))

	.dataa(!din_a[182]),
	.datab(!din_b[186]),
	.datac(!din_a[183]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_341 ),
	.sharein(Xd_0__inst_mult_15_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_468 ),
	.cout(Xd_0__inst_mult_15_469 ),
	.shareout(Xd_0__inst_mult_15_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_143 (
// Equation(s):
// Xd_0__inst_mult_15_473  = CARRY(( GND ) + ( Xd_0__inst_i29_55  ) + ( Xd_0__inst_i29_54  ))
// Xd_0__inst_mult_15_474  = SHARE((din_a[180] & din_b[188]))

	.dataa(!din_a[180]),
	.datab(!din_b[188]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_54 ),
	.sharein(Xd_0__inst_i29_55 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_473 ),
	.shareout(Xd_0__inst_mult_15_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_129 (
// Equation(s):
// Xd_0__inst_mult_10_428  = SUM(( (din_a[126] & din_b[122]) ) + ( Xd_0__inst_mult_10_422  ) + ( Xd_0__inst_mult_10_421  ))
// Xd_0__inst_mult_10_429  = CARRY(( (din_a[126] & din_b[122]) ) + ( Xd_0__inst_mult_10_422  ) + ( Xd_0__inst_mult_10_421  ))
// Xd_0__inst_mult_10_430  = SHARE((din_a[128] & din_b[121]))

	.dataa(!din_a[126]),
	.datab(!din_b[122]),
	.datac(!din_a[128]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_421 ),
	.sharein(Xd_0__inst_mult_10_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_428 ),
	.cout(Xd_0__inst_mult_10_429 ),
	.shareout(Xd_0__inst_mult_10_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_130 (
// Equation(s):
// Xd_0__inst_mult_10_432  = SUM(( (!din_a[125] & (((din_a[124] & din_b[124])))) # (din_a[125] & (!din_b[123] $ (((!din_a[124]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_426  ) + ( Xd_0__inst_mult_10_425  ))
// Xd_0__inst_mult_10_433  = CARRY(( (!din_a[125] & (((din_a[124] & din_b[124])))) # (din_a[125] & (!din_b[123] $ (((!din_a[124]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_426  ) + ( Xd_0__inst_mult_10_425  ))
// Xd_0__inst_mult_10_434  = SHARE((din_a[125] & (din_b[123] & (din_a[124] & din_b[124]))))

	.dataa(!din_a[125]),
	.datab(!din_b[123]),
	.datac(!din_a[124]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_425 ),
	.sharein(Xd_0__inst_mult_10_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_432 ),
	.cout(Xd_0__inst_mult_10_433 ),
	.shareout(Xd_0__inst_mult_10_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_131 (
// Equation(s):
// Xd_0__inst_mult_10_436  = SUM(( (!din_a[122] & (((din_a[123] & din_b[125])))) # (din_a[122] & (!din_b[126] $ (((!din_a[123]) # (!din_b[125]))))) ) + ( Xd_0__inst_mult_10_314  ) + ( Xd_0__inst_mult_10_313  ))
// Xd_0__inst_mult_10_437  = CARRY(( (!din_a[122] & (((din_a[123] & din_b[125])))) # (din_a[122] & (!din_b[126] $ (((!din_a[123]) # (!din_b[125]))))) ) + ( Xd_0__inst_mult_10_314  ) + ( Xd_0__inst_mult_10_313  ))
// Xd_0__inst_mult_10_438  = SHARE((din_a[122] & (din_b[126] & (din_a[123] & din_b[125]))))

	.dataa(!din_a[122]),
	.datab(!din_b[126]),
	.datac(!din_a[123]),
	.datad(!din_b[125]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_313 ),
	.sharein(Xd_0__inst_mult_10_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_436 ),
	.cout(Xd_0__inst_mult_10_437 ),
	.shareout(Xd_0__inst_mult_10_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_132 (
// Equation(s):
// Xd_0__inst_mult_10_441  = CARRY(( GND ) + ( Xd_0__inst_mult_2_53  ) + ( Xd_0__inst_mult_2_52  ))
// Xd_0__inst_mult_10_442  = SHARE((din_a[120] & din_b[128]))

	.dataa(!din_a[120]),
	.datab(!din_b[128]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_52 ),
	.sharein(Xd_0__inst_mult_2_53 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_441 ),
	.shareout(Xd_0__inst_mult_10_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_133 (
// Equation(s):
// Xd_0__inst_mult_11_432  = SUM(( (din_a[138] & din_b[134]) ) + ( Xd_0__inst_mult_11_426  ) + ( Xd_0__inst_mult_11_425  ))
// Xd_0__inst_mult_11_433  = CARRY(( (din_a[138] & din_b[134]) ) + ( Xd_0__inst_mult_11_426  ) + ( Xd_0__inst_mult_11_425  ))
// Xd_0__inst_mult_11_434  = SHARE((din_a[140] & din_b[133]))

	.dataa(!din_a[138]),
	.datab(!din_b[134]),
	.datac(!din_a[140]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_425 ),
	.sharein(Xd_0__inst_mult_11_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_432 ),
	.cout(Xd_0__inst_mult_11_433 ),
	.shareout(Xd_0__inst_mult_11_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_134 (
// Equation(s):
// Xd_0__inst_mult_11_436  = SUM(( (!din_a[137] & (((din_a[136] & din_b[136])))) # (din_a[137] & (!din_b[135] $ (((!din_a[136]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_430  ) + ( Xd_0__inst_mult_11_429  ))
// Xd_0__inst_mult_11_437  = CARRY(( (!din_a[137] & (((din_a[136] & din_b[136])))) # (din_a[137] & (!din_b[135] $ (((!din_a[136]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_430  ) + ( Xd_0__inst_mult_11_429  ))
// Xd_0__inst_mult_11_438  = SHARE((din_a[137] & (din_b[135] & (din_a[136] & din_b[136]))))

	.dataa(!din_a[137]),
	.datab(!din_b[135]),
	.datac(!din_a[136]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_429 ),
	.sharein(Xd_0__inst_mult_11_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_436 ),
	.cout(Xd_0__inst_mult_11_437 ),
	.shareout(Xd_0__inst_mult_11_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_135 (
// Equation(s):
// Xd_0__inst_mult_11_440  = SUM(( (!din_a[134] & (((din_a[135] & din_b[137])))) # (din_a[134] & (!din_b[138] $ (((!din_a[135]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_11_318  ) + ( Xd_0__inst_mult_11_317  ))
// Xd_0__inst_mult_11_441  = CARRY(( (!din_a[134] & (((din_a[135] & din_b[137])))) # (din_a[134] & (!din_b[138] $ (((!din_a[135]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_11_318  ) + ( Xd_0__inst_mult_11_317  ))
// Xd_0__inst_mult_11_442  = SHARE((din_a[134] & (din_b[138] & (din_a[135] & din_b[137]))))

	.dataa(!din_a[134]),
	.datab(!din_b[138]),
	.datac(!din_a[135]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_317 ),
	.sharein(Xd_0__inst_mult_11_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_440 ),
	.cout(Xd_0__inst_mult_11_441 ),
	.shareout(Xd_0__inst_mult_11_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_136 (
// Equation(s):
// Xd_0__inst_mult_11_445  = CARRY(( GND ) + ( Xd_0__inst_mult_12_61  ) + ( Xd_0__inst_mult_12_60  ))
// Xd_0__inst_mult_11_446  = SHARE((din_a[132] & din_b[140]))

	.dataa(!din_a[132]),
	.datab(!din_b[140]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_60 ),
	.sharein(Xd_0__inst_mult_12_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_445 ),
	.shareout(Xd_0__inst_mult_11_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_133 (
// Equation(s):
// Xd_0__inst_mult_8_432  = SUM(( (din_a[102] & din_b[98]) ) + ( Xd_0__inst_mult_8_426  ) + ( Xd_0__inst_mult_8_425  ))
// Xd_0__inst_mult_8_433  = CARRY(( (din_a[102] & din_b[98]) ) + ( Xd_0__inst_mult_8_426  ) + ( Xd_0__inst_mult_8_425  ))
// Xd_0__inst_mult_8_434  = SHARE((din_a[104] & din_b[97]))

	.dataa(!din_a[102]),
	.datab(!din_b[98]),
	.datac(!din_a[104]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_425 ),
	.sharein(Xd_0__inst_mult_8_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_432 ),
	.cout(Xd_0__inst_mult_8_433 ),
	.shareout(Xd_0__inst_mult_8_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_134 (
// Equation(s):
// Xd_0__inst_mult_8_436  = SUM(( (!din_a[101] & (((din_a[100] & din_b[100])))) # (din_a[101] & (!din_b[99] $ (((!din_a[100]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_430  ) + ( Xd_0__inst_mult_8_429  ))
// Xd_0__inst_mult_8_437  = CARRY(( (!din_a[101] & (((din_a[100] & din_b[100])))) # (din_a[101] & (!din_b[99] $ (((!din_a[100]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_430  ) + ( Xd_0__inst_mult_8_429  ))
// Xd_0__inst_mult_8_438  = SHARE((din_a[101] & (din_b[99] & (din_a[100] & din_b[100]))))

	.dataa(!din_a[101]),
	.datab(!din_b[99]),
	.datac(!din_a[100]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_429 ),
	.sharein(Xd_0__inst_mult_8_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_436 ),
	.cout(Xd_0__inst_mult_8_437 ),
	.shareout(Xd_0__inst_mult_8_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_135 (
// Equation(s):
// Xd_0__inst_mult_8_440  = SUM(( (!din_a[98] & (((din_a[99] & din_b[101])))) # (din_a[98] & (!din_b[102] $ (((!din_a[99]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_8_318  ) + ( Xd_0__inst_mult_8_317  ))
// Xd_0__inst_mult_8_441  = CARRY(( (!din_a[98] & (((din_a[99] & din_b[101])))) # (din_a[98] & (!din_b[102] $ (((!din_a[99]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_8_318  ) + ( Xd_0__inst_mult_8_317  ))
// Xd_0__inst_mult_8_442  = SHARE((din_a[98] & (din_b[102] & (din_a[99] & din_b[101]))))

	.dataa(!din_a[98]),
	.datab(!din_b[102]),
	.datac(!din_a[99]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_317 ),
	.sharein(Xd_0__inst_mult_8_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_440 ),
	.cout(Xd_0__inst_mult_8_441 ),
	.shareout(Xd_0__inst_mult_8_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_136 (
// Equation(s):
// Xd_0__inst_mult_8_445  = CARRY(( GND ) + ( Xd_0__inst_mult_6_57  ) + ( Xd_0__inst_mult_6_56  ))
// Xd_0__inst_mult_8_446  = SHARE((din_a[96] & din_b[104]))

	.dataa(!din_a[96]),
	.datab(!din_b[104]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_56 ),
	.sharein(Xd_0__inst_mult_6_57 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_445 ),
	.shareout(Xd_0__inst_mult_8_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_129 (
// Equation(s):
// Xd_0__inst_mult_9_428  = SUM(( (din_a[114] & din_b[110]) ) + ( Xd_0__inst_mult_9_422  ) + ( Xd_0__inst_mult_9_421  ))
// Xd_0__inst_mult_9_429  = CARRY(( (din_a[114] & din_b[110]) ) + ( Xd_0__inst_mult_9_422  ) + ( Xd_0__inst_mult_9_421  ))
// Xd_0__inst_mult_9_430  = SHARE((din_a[116] & din_b[109]))

	.dataa(!din_a[114]),
	.datab(!din_b[110]),
	.datac(!din_a[116]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_421 ),
	.sharein(Xd_0__inst_mult_9_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_428 ),
	.cout(Xd_0__inst_mult_9_429 ),
	.shareout(Xd_0__inst_mult_9_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_130 (
// Equation(s):
// Xd_0__inst_mult_9_432  = SUM(( (!din_a[113] & (((din_a[112] & din_b[112])))) # (din_a[113] & (!din_b[111] $ (((!din_a[112]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_426  ) + ( Xd_0__inst_mult_9_425  ))
// Xd_0__inst_mult_9_433  = CARRY(( (!din_a[113] & (((din_a[112] & din_b[112])))) # (din_a[113] & (!din_b[111] $ (((!din_a[112]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_426  ) + ( Xd_0__inst_mult_9_425  ))
// Xd_0__inst_mult_9_434  = SHARE((din_a[113] & (din_b[111] & (din_a[112] & din_b[112]))))

	.dataa(!din_a[113]),
	.datab(!din_b[111]),
	.datac(!din_a[112]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_425 ),
	.sharein(Xd_0__inst_mult_9_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_432 ),
	.cout(Xd_0__inst_mult_9_433 ),
	.shareout(Xd_0__inst_mult_9_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_63 (
// Equation(s):
// Xd_0__inst_mult_9_63_sumout  = SUM(( (din_a[116] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_64  = CARRY(( (din_a[116] & din_b[108]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_65  = SHARE(GND)

	.dataa(!din_a[116]),
	.datab(!din_b[108]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_9_63_sumout ),
	.cout(Xd_0__inst_mult_9_64 ),
	.shareout(Xd_0__inst_mult_9_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_131 (
// Equation(s):
// Xd_0__inst_mult_9_436  = SUM(( (!din_a[110] & (((din_a[111] & din_b[113])))) # (din_a[110] & (!din_b[114] $ (((!din_a[111]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_9_314  ) + ( Xd_0__inst_mult_9_313  ))
// Xd_0__inst_mult_9_437  = CARRY(( (!din_a[110] & (((din_a[111] & din_b[113])))) # (din_a[110] & (!din_b[114] $ (((!din_a[111]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_9_314  ) + ( Xd_0__inst_mult_9_313  ))
// Xd_0__inst_mult_9_438  = SHARE((din_a[110] & (din_b[114] & (din_a[111] & din_b[113]))))

	.dataa(!din_a[110]),
	.datab(!din_b[114]),
	.datac(!din_a[111]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_313 ),
	.sharein(Xd_0__inst_mult_9_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_436 ),
	.cout(Xd_0__inst_mult_9_437 ),
	.shareout(Xd_0__inst_mult_9_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_132 (
// Equation(s):
// Xd_0__inst_mult_9_441  = CARRY(( GND ) + ( Xd_0__inst_mult_0_53  ) + ( Xd_0__inst_mult_0_52  ))
// Xd_0__inst_mult_9_442  = SHARE((din_a[108] & din_b[116]))

	.dataa(!din_a[108]),
	.datab(!din_b[116]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_52 ),
	.sharein(Xd_0__inst_mult_0_53 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_441 ),
	.shareout(Xd_0__inst_mult_9_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_129 (
// Equation(s):
// Xd_0__inst_mult_6_428  = SUM(( (din_a[78] & din_b[74]) ) + ( Xd_0__inst_mult_6_422  ) + ( Xd_0__inst_mult_6_421  ))
// Xd_0__inst_mult_6_429  = CARRY(( (din_a[78] & din_b[74]) ) + ( Xd_0__inst_mult_6_422  ) + ( Xd_0__inst_mult_6_421  ))
// Xd_0__inst_mult_6_430  = SHARE((din_a[80] & din_b[73]))

	.dataa(!din_a[78]),
	.datab(!din_b[74]),
	.datac(!din_a[80]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_421 ),
	.sharein(Xd_0__inst_mult_6_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_428 ),
	.cout(Xd_0__inst_mult_6_429 ),
	.shareout(Xd_0__inst_mult_6_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_130 (
// Equation(s):
// Xd_0__inst_mult_6_432  = SUM(( (!din_a[77] & (((din_a[76] & din_b[76])))) # (din_a[77] & (!din_b[75] $ (((!din_a[76]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_426  ) + ( Xd_0__inst_mult_6_425  ))
// Xd_0__inst_mult_6_433  = CARRY(( (!din_a[77] & (((din_a[76] & din_b[76])))) # (din_a[77] & (!din_b[75] $ (((!din_a[76]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_426  ) + ( Xd_0__inst_mult_6_425  ))
// Xd_0__inst_mult_6_434  = SHARE((din_a[77] & (din_b[75] & (din_a[76] & din_b[76]))))

	.dataa(!din_a[77]),
	.datab(!din_b[75]),
	.datac(!din_a[76]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_425 ),
	.sharein(Xd_0__inst_mult_6_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_432 ),
	.cout(Xd_0__inst_mult_6_433 ),
	.shareout(Xd_0__inst_mult_6_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_131 (
// Equation(s):
// Xd_0__inst_mult_6_436  = SUM(( (!din_a[74] & (((din_a[75] & din_b[77])))) # (din_a[74] & (!din_b[78] $ (((!din_a[75]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_314  ) + ( Xd_0__inst_mult_6_313  ))
// Xd_0__inst_mult_6_437  = CARRY(( (!din_a[74] & (((din_a[75] & din_b[77])))) # (din_a[74] & (!din_b[78] $ (((!din_a[75]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_314  ) + ( Xd_0__inst_mult_6_313  ))
// Xd_0__inst_mult_6_438  = SHARE((din_a[74] & (din_b[78] & (din_a[75] & din_b[77]))))

	.dataa(!din_a[74]),
	.datab(!din_b[78]),
	.datac(!din_a[75]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_313 ),
	.sharein(Xd_0__inst_mult_6_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_436 ),
	.cout(Xd_0__inst_mult_6_437 ),
	.shareout(Xd_0__inst_mult_6_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_132 (
// Equation(s):
// Xd_0__inst_mult_6_441  = CARRY(( GND ) + ( Xd_0__inst_mult_2_49  ) + ( Xd_0__inst_mult_2_48  ))
// Xd_0__inst_mult_6_442  = SHARE((din_a[72] & din_b[80]))

	.dataa(!din_a[72]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_48 ),
	.sharein(Xd_0__inst_mult_2_49 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_441 ),
	.shareout(Xd_0__inst_mult_6_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_125 (
// Equation(s):
// Xd_0__inst_mult_7_412  = SUM(( (din_a[90] & din_b[86]) ) + ( Xd_0__inst_mult_7_406  ) + ( Xd_0__inst_mult_7_405  ))
// Xd_0__inst_mult_7_413  = CARRY(( (din_a[90] & din_b[86]) ) + ( Xd_0__inst_mult_7_406  ) + ( Xd_0__inst_mult_7_405  ))
// Xd_0__inst_mult_7_414  = SHARE((din_a[92] & din_b[85]))

	.dataa(!din_a[90]),
	.datab(!din_b[86]),
	.datac(!din_a[92]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_405 ),
	.sharein(Xd_0__inst_mult_7_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_412 ),
	.cout(Xd_0__inst_mult_7_413 ),
	.shareout(Xd_0__inst_mult_7_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_126 (
// Equation(s):
// Xd_0__inst_mult_7_416  = SUM(( (!din_a[89] & (((din_a[88] & din_b[88])))) # (din_a[89] & (!din_b[87] $ (((!din_a[88]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_410  ) + ( Xd_0__inst_mult_7_409  ))
// Xd_0__inst_mult_7_417  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[88])))) # (din_a[89] & (!din_b[87] $ (((!din_a[88]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_410  ) + ( Xd_0__inst_mult_7_409  ))
// Xd_0__inst_mult_7_418  = SHARE((din_a[89] & (din_b[87] & (din_a[88] & din_b[88]))))

	.dataa(!din_a[89]),
	.datab(!din_b[87]),
	.datac(!din_a[88]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_409 ),
	.sharein(Xd_0__inst_mult_7_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_416 ),
	.cout(Xd_0__inst_mult_7_417 ),
	.shareout(Xd_0__inst_mult_7_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_59 (
// Equation(s):
// Xd_0__inst_mult_7_59_sumout  = SUM(( (din_a[92] & din_b[84]) ) + ( Xd_0__inst_mult_4_65  ) + ( Xd_0__inst_mult_4_64  ))
// Xd_0__inst_mult_7_60  = CARRY(( (din_a[92] & din_b[84]) ) + ( Xd_0__inst_mult_4_65  ) + ( Xd_0__inst_mult_4_64  ))
// Xd_0__inst_mult_7_61  = SHARE(GND)

	.dataa(!din_a[92]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_64 ),
	.sharein(Xd_0__inst_mult_4_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_59_sumout ),
	.cout(Xd_0__inst_mult_7_60 ),
	.shareout(Xd_0__inst_mult_7_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_127 (
// Equation(s):
// Xd_0__inst_mult_7_420  = SUM(( (!din_a[86] & (((din_a[87] & din_b[89])))) # (din_a[86] & (!din_b[90] $ (((!din_a[87]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_290  ) + ( Xd_0__inst_mult_7_289  ))
// Xd_0__inst_mult_7_421  = CARRY(( (!din_a[86] & (((din_a[87] & din_b[89])))) # (din_a[86] & (!din_b[90] $ (((!din_a[87]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_290  ) + ( Xd_0__inst_mult_7_289  ))
// Xd_0__inst_mult_7_422  = SHARE((din_a[86] & (din_b[90] & (din_a[87] & din_b[89]))))

	.dataa(!din_a[86]),
	.datab(!din_b[90]),
	.datac(!din_a[87]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_289 ),
	.sharein(Xd_0__inst_mult_7_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_420 ),
	.cout(Xd_0__inst_mult_7_421 ),
	.shareout(Xd_0__inst_mult_7_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_128 (
// Equation(s):
// Xd_0__inst_mult_7_425  = CARRY(( GND ) + ( Xd_0__inst_mult_12_57  ) + ( Xd_0__inst_mult_12_56  ))
// Xd_0__inst_mult_7_426  = SHARE((din_a[84] & din_b[92]))

	.dataa(!din_a[84]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_56 ),
	.sharein(Xd_0__inst_mult_12_57 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_425 ),
	.shareout(Xd_0__inst_mult_7_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_138 (
// Equation(s):
// Xd_0__inst_mult_4_452  = SUM(( (din_a[54] & din_b[50]) ) + ( Xd_0__inst_mult_4_446  ) + ( Xd_0__inst_mult_4_445  ))
// Xd_0__inst_mult_4_453  = CARRY(( (din_a[54] & din_b[50]) ) + ( Xd_0__inst_mult_4_446  ) + ( Xd_0__inst_mult_4_445  ))
// Xd_0__inst_mult_4_454  = SHARE((din_a[56] & din_b[49]))

	.dataa(!din_a[54]),
	.datab(!din_b[50]),
	.datac(!din_a[56]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_445 ),
	.sharein(Xd_0__inst_mult_4_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_452 ),
	.cout(Xd_0__inst_mult_4_453 ),
	.shareout(Xd_0__inst_mult_4_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_139 (
// Equation(s):
// Xd_0__inst_mult_4_456  = SUM(( (!din_a[53] & (((din_a[52] & din_b[52])))) # (din_a[53] & (!din_b[51] $ (((!din_a[52]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_450  ) + ( Xd_0__inst_mult_4_449  ))
// Xd_0__inst_mult_4_457  = CARRY(( (!din_a[53] & (((din_a[52] & din_b[52])))) # (din_a[53] & (!din_b[51] $ (((!din_a[52]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_450  ) + ( Xd_0__inst_mult_4_449  ))
// Xd_0__inst_mult_4_458  = SHARE((din_a[53] & (din_b[51] & (din_a[52] & din_b[52]))))

	.dataa(!din_a[53]),
	.datab(!din_b[51]),
	.datac(!din_a[52]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_449 ),
	.sharein(Xd_0__inst_mult_4_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_456 ),
	.cout(Xd_0__inst_mult_4_457 ),
	.shareout(Xd_0__inst_mult_4_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_63 (
// Equation(s):
// Xd_0__inst_mult_4_63_sumout  = SUM(( (din_a[56] & din_b[48]) ) + ( Xd_0__inst_mult_5_65  ) + ( Xd_0__inst_mult_5_64  ))
// Xd_0__inst_mult_4_64  = CARRY(( (din_a[56] & din_b[48]) ) + ( Xd_0__inst_mult_5_65  ) + ( Xd_0__inst_mult_5_64  ))
// Xd_0__inst_mult_4_65  = SHARE(GND)

	.dataa(!din_a[56]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_64 ),
	.sharein(Xd_0__inst_mult_5_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_63_sumout ),
	.cout(Xd_0__inst_mult_4_64 ),
	.shareout(Xd_0__inst_mult_4_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_140 (
// Equation(s):
// Xd_0__inst_mult_4_460  = SUM(( (!din_a[50] & (((din_a[51] & din_b[53])))) # (din_a[50] & (!din_b[54] $ (((!din_a[51]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_326  ) + ( Xd_0__inst_mult_4_325  ))
// Xd_0__inst_mult_4_461  = CARRY(( (!din_a[50] & (((din_a[51] & din_b[53])))) # (din_a[50] & (!din_b[54] $ (((!din_a[51]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_326  ) + ( Xd_0__inst_mult_4_325  ))
// Xd_0__inst_mult_4_462  = SHARE((din_a[50] & (din_b[54] & (din_a[51] & din_b[53]))))

	.dataa(!din_a[50]),
	.datab(!din_b[54]),
	.datac(!din_a[51]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_325 ),
	.sharein(Xd_0__inst_mult_4_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_460 ),
	.cout(Xd_0__inst_mult_4_461 ),
	.shareout(Xd_0__inst_mult_4_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_141 (
// Equation(s):
// Xd_0__inst_mult_4_465  = CARRY(( GND ) + ( Xd_0__inst_mult_6_53  ) + ( Xd_0__inst_mult_6_52  ))
// Xd_0__inst_mult_4_466  = SHARE((din_a[48] & din_b[56]))

	.dataa(!din_a[48]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_52 ),
	.sharein(Xd_0__inst_mult_6_53 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_465 ),
	.shareout(Xd_0__inst_mult_4_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_125 (
// Equation(s):
// Xd_0__inst_mult_5_412  = SUM(( (din_a[66] & din_b[62]) ) + ( Xd_0__inst_mult_5_406  ) + ( Xd_0__inst_mult_5_405  ))
// Xd_0__inst_mult_5_413  = CARRY(( (din_a[66] & din_b[62]) ) + ( Xd_0__inst_mult_5_406  ) + ( Xd_0__inst_mult_5_405  ))
// Xd_0__inst_mult_5_414  = SHARE((din_a[68] & din_b[61]))

	.dataa(!din_a[66]),
	.datab(!din_b[62]),
	.datac(!din_a[68]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_405 ),
	.sharein(Xd_0__inst_mult_5_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_412 ),
	.cout(Xd_0__inst_mult_5_413 ),
	.shareout(Xd_0__inst_mult_5_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_126 (
// Equation(s):
// Xd_0__inst_mult_5_416  = SUM(( (!din_a[65] & (((din_a[64] & din_b[64])))) # (din_a[65] & (!din_b[63] $ (((!din_a[64]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_410  ) + ( Xd_0__inst_mult_5_409  ))
// Xd_0__inst_mult_5_417  = CARRY(( (!din_a[65] & (((din_a[64] & din_b[64])))) # (din_a[65] & (!din_b[63] $ (((!din_a[64]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_410  ) + ( Xd_0__inst_mult_5_409  ))
// Xd_0__inst_mult_5_418  = SHARE((din_a[65] & (din_b[63] & (din_a[64] & din_b[64]))))

	.dataa(!din_a[65]),
	.datab(!din_b[63]),
	.datac(!din_a[64]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_409 ),
	.sharein(Xd_0__inst_mult_5_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_416 ),
	.cout(Xd_0__inst_mult_5_417 ),
	.shareout(Xd_0__inst_mult_5_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_63 (
// Equation(s):
// Xd_0__inst_mult_5_63_sumout  = SUM(( (din_a[68] & din_b[60]) ) + ( Xd_0__inst_mult_2_65  ) + ( Xd_0__inst_mult_2_64  ))
// Xd_0__inst_mult_5_64  = CARRY(( (din_a[68] & din_b[60]) ) + ( Xd_0__inst_mult_2_65  ) + ( Xd_0__inst_mult_2_64  ))
// Xd_0__inst_mult_5_65  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_64 ),
	.sharein(Xd_0__inst_mult_2_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_63_sumout ),
	.cout(Xd_0__inst_mult_5_64 ),
	.shareout(Xd_0__inst_mult_5_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_127 (
// Equation(s):
// Xd_0__inst_mult_5_420  = SUM(( (!din_a[62] & (((din_a[63] & din_b[65])))) # (din_a[62] & (!din_b[66] $ (((!din_a[63]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_290  ) + ( Xd_0__inst_mult_5_289  ))
// Xd_0__inst_mult_5_421  = CARRY(( (!din_a[62] & (((din_a[63] & din_b[65])))) # (din_a[62] & (!din_b[66] $ (((!din_a[63]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_290  ) + ( Xd_0__inst_mult_5_289  ))
// Xd_0__inst_mult_5_422  = SHARE((din_a[62] & (din_b[66] & (din_a[63] & din_b[65]))))

	.dataa(!din_a[62]),
	.datab(!din_b[66]),
	.datac(!din_a[63]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_289 ),
	.sharein(Xd_0__inst_mult_5_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_420 ),
	.cout(Xd_0__inst_mult_5_421 ),
	.shareout(Xd_0__inst_mult_5_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_128 (
// Equation(s):
// Xd_0__inst_mult_5_425  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_426  = SHARE((din_a[60] & din_b[68]))

	.dataa(!din_a[60]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_425 ),
	.shareout(Xd_0__inst_mult_5_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_129 (
// Equation(s):
// Xd_0__inst_mult_2_416  = SUM(( (din_a[30] & din_b[26]) ) + ( Xd_0__inst_mult_2_410  ) + ( Xd_0__inst_mult_2_409  ))
// Xd_0__inst_mult_2_417  = CARRY(( (din_a[30] & din_b[26]) ) + ( Xd_0__inst_mult_2_410  ) + ( Xd_0__inst_mult_2_409  ))
// Xd_0__inst_mult_2_418  = SHARE((din_a[32] & din_b[25]))

	.dataa(!din_a[30]),
	.datab(!din_b[26]),
	.datac(!din_a[32]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_409 ),
	.sharein(Xd_0__inst_mult_2_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_416 ),
	.cout(Xd_0__inst_mult_2_417 ),
	.shareout(Xd_0__inst_mult_2_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_130 (
// Equation(s):
// Xd_0__inst_mult_2_420  = SUM(( (!din_a[29] & (((din_a[28] & din_b[28])))) # (din_a[29] & (!din_b[27] $ (((!din_a[28]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_414  ) + ( Xd_0__inst_mult_2_413  ))
// Xd_0__inst_mult_2_421  = CARRY(( (!din_a[29] & (((din_a[28] & din_b[28])))) # (din_a[29] & (!din_b[27] $ (((!din_a[28]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_414  ) + ( Xd_0__inst_mult_2_413  ))
// Xd_0__inst_mult_2_422  = SHARE((din_a[29] & (din_b[27] & (din_a[28] & din_b[28]))))

	.dataa(!din_a[29]),
	.datab(!din_b[27]),
	.datac(!din_a[28]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_413 ),
	.sharein(Xd_0__inst_mult_2_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_420 ),
	.cout(Xd_0__inst_mult_2_421 ),
	.shareout(Xd_0__inst_mult_2_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_63 (
// Equation(s):
// Xd_0__inst_mult_2_63_sumout  = SUM(( (din_a[32] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_64  = CARRY(( (din_a[32] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_65  = SHARE(GND)

	.dataa(!din_a[32]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_63_sumout ),
	.cout(Xd_0__inst_mult_2_64 ),
	.shareout(Xd_0__inst_mult_2_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_131 (
// Equation(s):
// Xd_0__inst_mult_2_424  = SUM(( (!din_a[26] & (((din_a[27] & din_b[29])))) # (din_a[26] & (!din_b[30] $ (((!din_a[27]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_294  ) + ( Xd_0__inst_mult_2_293  ))
// Xd_0__inst_mult_2_425  = CARRY(( (!din_a[26] & (((din_a[27] & din_b[29])))) # (din_a[26] & (!din_b[30] $ (((!din_a[27]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_294  ) + ( Xd_0__inst_mult_2_293  ))
// Xd_0__inst_mult_2_426  = SHARE((din_a[26] & (din_b[30] & (din_a[27] & din_b[29]))))

	.dataa(!din_a[26]),
	.datab(!din_b[30]),
	.datac(!din_a[27]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_293 ),
	.sharein(Xd_0__inst_mult_2_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_424 ),
	.cout(Xd_0__inst_mult_2_425 ),
	.shareout(Xd_0__inst_mult_2_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_132 (
// Equation(s):
// Xd_0__inst_mult_2_429  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_430  = SHARE((din_a[24] & din_b[32]))

	.dataa(!din_a[24]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_429 ),
	.shareout(Xd_0__inst_mult_2_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_125 (
// Equation(s):
// Xd_0__inst_mult_3_412  = SUM(( (din_a[42] & din_b[38]) ) + ( Xd_0__inst_mult_3_406  ) + ( Xd_0__inst_mult_3_405  ))
// Xd_0__inst_mult_3_413  = CARRY(( (din_a[42] & din_b[38]) ) + ( Xd_0__inst_mult_3_406  ) + ( Xd_0__inst_mult_3_405  ))
// Xd_0__inst_mult_3_414  = SHARE((din_a[44] & din_b[37]))

	.dataa(!din_a[42]),
	.datab(!din_b[38]),
	.datac(!din_a[44]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_405 ),
	.sharein(Xd_0__inst_mult_3_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_412 ),
	.cout(Xd_0__inst_mult_3_413 ),
	.shareout(Xd_0__inst_mult_3_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_126 (
// Equation(s):
// Xd_0__inst_mult_3_416  = SUM(( (!din_a[41] & (((din_a[40] & din_b[40])))) # (din_a[41] & (!din_b[39] $ (((!din_a[40]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_410  ) + ( Xd_0__inst_mult_3_409  ))
// Xd_0__inst_mult_3_417  = CARRY(( (!din_a[41] & (((din_a[40] & din_b[40])))) # (din_a[41] & (!din_b[39] $ (((!din_a[40]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_410  ) + ( Xd_0__inst_mult_3_409  ))
// Xd_0__inst_mult_3_418  = SHARE((din_a[41] & (din_b[39] & (din_a[40] & din_b[40]))))

	.dataa(!din_a[41]),
	.datab(!din_b[39]),
	.datac(!din_a[40]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_409 ),
	.sharein(Xd_0__inst_mult_3_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_416 ),
	.cout(Xd_0__inst_mult_3_417 ),
	.shareout(Xd_0__inst_mult_3_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_127 (
// Equation(s):
// Xd_0__inst_mult_3_420  = SUM(( (!din_a[38] & (((din_a[39] & din_b[41])))) # (din_a[38] & (!din_b[42] $ (((!din_a[39]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_290  ) + ( Xd_0__inst_mult_3_289  ))
// Xd_0__inst_mult_3_421  = CARRY(( (!din_a[38] & (((din_a[39] & din_b[41])))) # (din_a[38] & (!din_b[42] $ (((!din_a[39]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_290  ) + ( Xd_0__inst_mult_3_289  ))
// Xd_0__inst_mult_3_422  = SHARE((din_a[38] & (din_b[42] & (din_a[39] & din_b[41]))))

	.dataa(!din_a[38]),
	.datab(!din_b[42]),
	.datac(!din_a[39]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_289 ),
	.sharein(Xd_0__inst_mult_3_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_420 ),
	.cout(Xd_0__inst_mult_3_421 ),
	.shareout(Xd_0__inst_mult_3_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_128 (
// Equation(s):
// Xd_0__inst_mult_3_425  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_426  = SHARE((din_a[36] & din_b[44]))

	.dataa(!din_a[36]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_425 ),
	.shareout(Xd_0__inst_mult_3_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_129 (
// Equation(s):
// Xd_0__inst_mult_0_416  = SUM(( (din_a[6] & din_b[2]) ) + ( Xd_0__inst_mult_0_410  ) + ( Xd_0__inst_mult_0_409  ))
// Xd_0__inst_mult_0_417  = CARRY(( (din_a[6] & din_b[2]) ) + ( Xd_0__inst_mult_0_410  ) + ( Xd_0__inst_mult_0_409  ))
// Xd_0__inst_mult_0_418  = SHARE((din_a[8] & din_b[1]))

	.dataa(!din_a[6]),
	.datab(!din_b[2]),
	.datac(!din_a[8]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_409 ),
	.sharein(Xd_0__inst_mult_0_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_416 ),
	.cout(Xd_0__inst_mult_0_417 ),
	.shareout(Xd_0__inst_mult_0_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_130 (
// Equation(s):
// Xd_0__inst_mult_0_420  = SUM(( (!din_a[5] & (((din_a[4] & din_b[4])))) # (din_a[5] & (!din_b[3] $ (((!din_a[4]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_414  ) + ( Xd_0__inst_mult_0_413  ))
// Xd_0__inst_mult_0_421  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[4])))) # (din_a[5] & (!din_b[3] $ (((!din_a[4]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_414  ) + ( Xd_0__inst_mult_0_413  ))
// Xd_0__inst_mult_0_422  = SHARE((din_a[5] & (din_b[3] & (din_a[4] & din_b[4]))))

	.dataa(!din_a[5]),
	.datab(!din_b[3]),
	.datac(!din_a[4]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_413 ),
	.sharein(Xd_0__inst_mult_0_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_420 ),
	.cout(Xd_0__inst_mult_0_421 ),
	.shareout(Xd_0__inst_mult_0_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_63 (
// Equation(s):
// Xd_0__inst_mult_0_63_sumout  = SUM(( (din_a[8] & din_b[0]) ) + ( Xd_0__inst_mult_1_69  ) + ( Xd_0__inst_mult_1_68  ))
// Xd_0__inst_mult_0_64  = CARRY(( (din_a[8] & din_b[0]) ) + ( Xd_0__inst_mult_1_69  ) + ( Xd_0__inst_mult_1_68  ))
// Xd_0__inst_mult_0_65  = SHARE(GND)

	.dataa(!din_a[8]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_68 ),
	.sharein(Xd_0__inst_mult_1_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_63_sumout ),
	.cout(Xd_0__inst_mult_0_64 ),
	.shareout(Xd_0__inst_mult_0_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_131 (
// Equation(s):
// Xd_0__inst_mult_0_424  = SUM(( (!din_a[2] & (((din_a[3] & din_b[5])))) # (din_a[2] & (!din_b[6] $ (((!din_a[3]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_294  ) + ( Xd_0__inst_mult_0_293  ))
// Xd_0__inst_mult_0_425  = CARRY(( (!din_a[2] & (((din_a[3] & din_b[5])))) # (din_a[2] & (!din_b[6] $ (((!din_a[3]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_294  ) + ( Xd_0__inst_mult_0_293  ))
// Xd_0__inst_mult_0_426  = SHARE((din_a[2] & (din_b[6] & (din_a[3] & din_b[5]))))

	.dataa(!din_a[2]),
	.datab(!din_b[6]),
	.datac(!din_a[3]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_293 ),
	.sharein(Xd_0__inst_mult_0_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_424 ),
	.cout(Xd_0__inst_mult_0_425 ),
	.shareout(Xd_0__inst_mult_0_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_132 (
// Equation(s):
// Xd_0__inst_mult_0_429  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_430  = SHARE((din_a[0] & din_b[8]))

	.dataa(!din_a[0]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_429 ),
	.shareout(Xd_0__inst_mult_0_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_129 (
// Equation(s):
// Xd_0__inst_mult_1_416  = SUM(( (din_a[18] & din_b[14]) ) + ( Xd_0__inst_mult_1_410  ) + ( Xd_0__inst_mult_1_409  ))
// Xd_0__inst_mult_1_417  = CARRY(( (din_a[18] & din_b[14]) ) + ( Xd_0__inst_mult_1_410  ) + ( Xd_0__inst_mult_1_409  ))
// Xd_0__inst_mult_1_418  = SHARE((din_a[20] & din_b[13]))

	.dataa(!din_a[18]),
	.datab(!din_b[14]),
	.datac(!din_a[20]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_409 ),
	.sharein(Xd_0__inst_mult_1_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_416 ),
	.cout(Xd_0__inst_mult_1_417 ),
	.shareout(Xd_0__inst_mult_1_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_130 (
// Equation(s):
// Xd_0__inst_mult_1_420  = SUM(( (!din_a[17] & (((din_a[16] & din_b[16])))) # (din_a[17] & (!din_b[15] $ (((!din_a[16]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_414  ) + ( Xd_0__inst_mult_1_413  ))
// Xd_0__inst_mult_1_421  = CARRY(( (!din_a[17] & (((din_a[16] & din_b[16])))) # (din_a[17] & (!din_b[15] $ (((!din_a[16]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_414  ) + ( Xd_0__inst_mult_1_413  ))
// Xd_0__inst_mult_1_422  = SHARE((din_a[17] & (din_b[15] & (din_a[16] & din_b[16]))))

	.dataa(!din_a[17]),
	.datab(!din_b[15]),
	.datac(!din_a[16]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_413 ),
	.sharein(Xd_0__inst_mult_1_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_420 ),
	.cout(Xd_0__inst_mult_1_421 ),
	.shareout(Xd_0__inst_mult_1_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_67 (
// Equation(s):
// Xd_0__inst_mult_1_67_sumout  = SUM(( (din_a[20] & din_b[12]) ) + ( Xd_0__inst_mult_14_69  ) + ( Xd_0__inst_mult_14_68  ))
// Xd_0__inst_mult_1_68  = CARRY(( (din_a[20] & din_b[12]) ) + ( Xd_0__inst_mult_14_69  ) + ( Xd_0__inst_mult_14_68  ))
// Xd_0__inst_mult_1_69  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_68 ),
	.sharein(Xd_0__inst_mult_14_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_67_sumout ),
	.cout(Xd_0__inst_mult_1_68 ),
	.shareout(Xd_0__inst_mult_1_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_131 (
// Equation(s):
// Xd_0__inst_mult_1_424  = SUM(( (!din_a[14] & (((din_a[15] & din_b[17])))) # (din_a[14] & (!din_b[18] $ (((!din_a[15]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_294  ) + ( Xd_0__inst_mult_1_293  ))
// Xd_0__inst_mult_1_425  = CARRY(( (!din_a[14] & (((din_a[15] & din_b[17])))) # (din_a[14] & (!din_b[18] $ (((!din_a[15]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_294  ) + ( Xd_0__inst_mult_1_293  ))
// Xd_0__inst_mult_1_426  = SHARE((din_a[14] & (din_b[18] & (din_a[15] & din_b[17]))))

	.dataa(!din_a[14]),
	.datab(!din_b[18]),
	.datac(!din_a[15]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_293 ),
	.sharein(Xd_0__inst_mult_1_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_424 ),
	.cout(Xd_0__inst_mult_1_425 ),
	.shareout(Xd_0__inst_mult_1_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_132 (
// Equation(s):
// Xd_0__inst_mult_1_429  = CARRY(( GND ) + ( Xd_0__inst_mult_0_41  ) + ( Xd_0__inst_mult_0_40  ))
// Xd_0__inst_mult_1_430  = SHARE((din_a[12] & din_b[20]))

	.dataa(!din_a[12]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_40 ),
	.sharein(Xd_0__inst_mult_0_41 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_429 ),
	.shareout(Xd_0__inst_mult_1_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_140 (
// Equation(s):
// Xd_0__inst_mult_12_472  = SUM(( (din_a[151] & din_b[146]) ) + ( Xd_0__inst_mult_12_458  ) + ( Xd_0__inst_mult_12_457  ))
// Xd_0__inst_mult_12_473  = CARRY(( (din_a[151] & din_b[146]) ) + ( Xd_0__inst_mult_12_458  ) + ( Xd_0__inst_mult_12_457  ))
// Xd_0__inst_mult_12_474  = SHARE((din_a[153] & din_b[145]))

	.dataa(!din_a[151]),
	.datab(!din_b[146]),
	.datac(!din_a[153]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_457 ),
	.sharein(Xd_0__inst_mult_12_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_472 ),
	.cout(Xd_0__inst_mult_12_473 ),
	.shareout(Xd_0__inst_mult_12_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_141 (
// Equation(s):
// Xd_0__inst_mult_12_476  = SUM(( (!din_a[150] & (((din_a[149] & din_b[148])))) # (din_a[150] & (!din_b[147] $ (((!din_a[149]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_462  ) + ( Xd_0__inst_mult_12_461  ))
// Xd_0__inst_mult_12_477  = CARRY(( (!din_a[150] & (((din_a[149] & din_b[148])))) # (din_a[150] & (!din_b[147] $ (((!din_a[149]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_462  ) + ( Xd_0__inst_mult_12_461  ))
// Xd_0__inst_mult_12_478  = SHARE((din_a[150] & (din_b[147] & (din_a[149] & din_b[148]))))

	.dataa(!din_a[150]),
	.datab(!din_b[147]),
	.datac(!din_a[149]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_461 ),
	.sharein(Xd_0__inst_mult_12_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_476 ),
	.cout(Xd_0__inst_mult_12_477 ),
	.shareout(Xd_0__inst_mult_12_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_142 (
// Equation(s):
// Xd_0__inst_mult_12_480  = SUM(( (!din_a[147] & (((din_a[148] & din_b[149])))) # (din_a[147] & (!din_b[150] $ (((!din_a[148]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_12_466  ) + ( Xd_0__inst_mult_12_465  ))
// Xd_0__inst_mult_12_481  = CARRY(( (!din_a[147] & (((din_a[148] & din_b[149])))) # (din_a[147] & (!din_b[150] $ (((!din_a[148]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_12_466  ) + ( Xd_0__inst_mult_12_465  ))
// Xd_0__inst_mult_12_482  = SHARE((din_a[147] & (din_b[150] & (din_a[148] & din_b[149]))))

	.dataa(!din_a[147]),
	.datab(!din_b[150]),
	.datac(!din_a[148]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_465 ),
	.sharein(Xd_0__inst_mult_12_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_480 ),
	.cout(Xd_0__inst_mult_12_481 ),
	.shareout(Xd_0__inst_mult_12_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_143 (
// Equation(s):
// Xd_0__inst_mult_12_484  = SUM(( (din_a[144] & din_b[153]) ) + ( Xd_0__inst_mult_12_574  ) + ( Xd_0__inst_mult_12_573  ))
// Xd_0__inst_mult_12_485  = CARRY(( (din_a[144] & din_b[153]) ) + ( Xd_0__inst_mult_12_574  ) + ( Xd_0__inst_mult_12_573  ))
// Xd_0__inst_mult_12_486  = SHARE((din_a[144] & din_b[154]))

	.dataa(!din_a[144]),
	.datab(!din_b[153]),
	.datac(!din_b[154]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_573 ),
	.sharein(Xd_0__inst_mult_12_574 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_484 ),
	.cout(Xd_0__inst_mult_12_485 ),
	.shareout(Xd_0__inst_mult_12_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_137 (
// Equation(s):
// Xd_0__inst_mult_13_448  = SUM(( (din_a[163] & din_b[158]) ) + ( Xd_0__inst_mult_13_434  ) + ( Xd_0__inst_mult_13_433  ))
// Xd_0__inst_mult_13_449  = CARRY(( (din_a[163] & din_b[158]) ) + ( Xd_0__inst_mult_13_434  ) + ( Xd_0__inst_mult_13_433  ))
// Xd_0__inst_mult_13_450  = SHARE((din_a[165] & din_b[157]))

	.dataa(!din_a[163]),
	.datab(!din_b[158]),
	.datac(!din_a[165]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_433 ),
	.sharein(Xd_0__inst_mult_13_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_448 ),
	.cout(Xd_0__inst_mult_13_449 ),
	.shareout(Xd_0__inst_mult_13_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_138 (
// Equation(s):
// Xd_0__inst_mult_13_452  = SUM(( (!din_a[162] & (((din_a[161] & din_b[160])))) # (din_a[162] & (!din_b[159] $ (((!din_a[161]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_438  ) + ( Xd_0__inst_mult_13_437  ))
// Xd_0__inst_mult_13_453  = CARRY(( (!din_a[162] & (((din_a[161] & din_b[160])))) # (din_a[162] & (!din_b[159] $ (((!din_a[161]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_438  ) + ( Xd_0__inst_mult_13_437  ))
// Xd_0__inst_mult_13_454  = SHARE((din_a[162] & (din_b[159] & (din_a[161] & din_b[160]))))

	.dataa(!din_a[162]),
	.datab(!din_b[159]),
	.datac(!din_a[161]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_437 ),
	.sharein(Xd_0__inst_mult_13_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_452 ),
	.cout(Xd_0__inst_mult_13_453 ),
	.shareout(Xd_0__inst_mult_13_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_67 (
// Equation(s):
// Xd_0__inst_mult_13_67_sumout  = SUM(( (din_a[165] & din_b[156]) ) + ( Xd_0__inst_mult_10_65  ) + ( Xd_0__inst_mult_10_64  ))
// Xd_0__inst_mult_13_68  = CARRY(( (din_a[165] & din_b[156]) ) + ( Xd_0__inst_mult_10_65  ) + ( Xd_0__inst_mult_10_64  ))
// Xd_0__inst_mult_13_69  = SHARE(GND)

	.dataa(!din_a[165]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_64 ),
	.sharein(Xd_0__inst_mult_10_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_67_sumout ),
	.cout(Xd_0__inst_mult_13_68 ),
	.shareout(Xd_0__inst_mult_13_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_139 (
// Equation(s):
// Xd_0__inst_mult_13_456  = SUM(( (!din_a[159] & (((din_a[160] & din_b[161])))) # (din_a[159] & (!din_b[162] $ (((!din_a[160]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_13_442  ) + ( Xd_0__inst_mult_13_441  ))
// Xd_0__inst_mult_13_457  = CARRY(( (!din_a[159] & (((din_a[160] & din_b[161])))) # (din_a[159] & (!din_b[162] $ (((!din_a[160]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_13_442  ) + ( Xd_0__inst_mult_13_441  ))
// Xd_0__inst_mult_13_458  = SHARE((din_a[159] & (din_b[162] & (din_a[160] & din_b[161]))))

	.dataa(!din_a[159]),
	.datab(!din_b[162]),
	.datac(!din_a[160]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_441 ),
	.sharein(Xd_0__inst_mult_13_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_456 ),
	.cout(Xd_0__inst_mult_13_457 ),
	.shareout(Xd_0__inst_mult_13_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_140 (
// Equation(s):
// Xd_0__inst_mult_13_460  = SUM(( (din_a[156] & din_b[165]) ) + ( Xd_0__inst_mult_13_582  ) + ( Xd_0__inst_mult_13_581  ))
// Xd_0__inst_mult_13_461  = CARRY(( (din_a[156] & din_b[165]) ) + ( Xd_0__inst_mult_13_582  ) + ( Xd_0__inst_mult_13_581  ))
// Xd_0__inst_mult_13_462  = SHARE((din_a[156] & din_b[166]))

	.dataa(!din_a[156]),
	.datab(!din_b[165]),
	.datac(!din_b[166]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_581 ),
	.sharein(Xd_0__inst_mult_13_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_460 ),
	.cout(Xd_0__inst_mult_13_461 ),
	.shareout(Xd_0__inst_mult_13_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_141 (
// Equation(s):
// Xd_0__inst_mult_14_464  = SUM(( (din_a[175] & din_b[170]) ) + ( Xd_0__inst_mult_14_450  ) + ( Xd_0__inst_mult_14_449  ))
// Xd_0__inst_mult_14_465  = CARRY(( (din_a[175] & din_b[170]) ) + ( Xd_0__inst_mult_14_450  ) + ( Xd_0__inst_mult_14_449  ))
// Xd_0__inst_mult_14_466  = SHARE((din_a[177] & din_b[169]))

	.dataa(!din_a[175]),
	.datab(!din_b[170]),
	.datac(!din_a[177]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_449 ),
	.sharein(Xd_0__inst_mult_14_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_464 ),
	.cout(Xd_0__inst_mult_14_465 ),
	.shareout(Xd_0__inst_mult_14_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_142 (
// Equation(s):
// Xd_0__inst_mult_14_468  = SUM(( (!din_a[174] & (((din_a[173] & din_b[172])))) # (din_a[174] & (!din_b[171] $ (((!din_a[173]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_454  ) + ( Xd_0__inst_mult_14_453  ))
// Xd_0__inst_mult_14_469  = CARRY(( (!din_a[174] & (((din_a[173] & din_b[172])))) # (din_a[174] & (!din_b[171] $ (((!din_a[173]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_14_454  ) + ( Xd_0__inst_mult_14_453  ))
// Xd_0__inst_mult_14_470  = SHARE((din_a[174] & (din_b[171] & (din_a[173] & din_b[172]))))

	.dataa(!din_a[174]),
	.datab(!din_b[171]),
	.datac(!din_a[173]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_453 ),
	.sharein(Xd_0__inst_mult_14_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_468 ),
	.cout(Xd_0__inst_mult_14_469 ),
	.shareout(Xd_0__inst_mult_14_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_67 (
// Equation(s):
// Xd_0__inst_mult_14_67_sumout  = SUM(( (din_a[177] & din_b[168]) ) + ( Xd_0__inst_mult_9_65  ) + ( Xd_0__inst_mult_9_64  ))
// Xd_0__inst_mult_14_68  = CARRY(( (din_a[177] & din_b[168]) ) + ( Xd_0__inst_mult_9_65  ) + ( Xd_0__inst_mult_9_64  ))
// Xd_0__inst_mult_14_69  = SHARE(GND)

	.dataa(!din_a[177]),
	.datab(!din_b[168]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_64 ),
	.sharein(Xd_0__inst_mult_9_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_67_sumout ),
	.cout(Xd_0__inst_mult_14_68 ),
	.shareout(Xd_0__inst_mult_14_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_143 (
// Equation(s):
// Xd_0__inst_mult_14_472  = SUM(( (!din_a[171] & (((din_a[172] & din_b[173])))) # (din_a[171] & (!din_b[174] $ (((!din_a[172]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_14_458  ) + ( Xd_0__inst_mult_14_457  ))
// Xd_0__inst_mult_14_473  = CARRY(( (!din_a[171] & (((din_a[172] & din_b[173])))) # (din_a[171] & (!din_b[174] $ (((!din_a[172]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_14_458  ) + ( Xd_0__inst_mult_14_457  ))
// Xd_0__inst_mult_14_474  = SHARE((din_a[171] & (din_b[174] & (din_a[172] & din_b[173]))))

	.dataa(!din_a[171]),
	.datab(!din_b[174]),
	.datac(!din_a[172]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_457 ),
	.sharein(Xd_0__inst_mult_14_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_472 ),
	.cout(Xd_0__inst_mult_14_473 ),
	.shareout(Xd_0__inst_mult_14_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_144 (
// Equation(s):
// Xd_0__inst_mult_14_476  = SUM(( (din_a[168] & din_b[177]) ) + ( Xd_0__inst_mult_14_582  ) + ( Xd_0__inst_mult_14_581  ))
// Xd_0__inst_mult_14_477  = CARRY(( (din_a[168] & din_b[177]) ) + ( Xd_0__inst_mult_14_582  ) + ( Xd_0__inst_mult_14_581  ))
// Xd_0__inst_mult_14_478  = SHARE((din_a[168] & din_b[178]))

	.dataa(!din_a[168]),
	.datab(!din_b[177]),
	.datac(!din_b[178]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_581 ),
	.sharein(Xd_0__inst_mult_14_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_476 ),
	.cout(Xd_0__inst_mult_14_477 ),
	.shareout(Xd_0__inst_mult_14_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_144 (
// Equation(s):
// Xd_0__inst_mult_15_476  = SUM(( (din_a[187] & din_b[182]) ) + ( Xd_0__inst_mult_15_462  ) + ( Xd_0__inst_mult_15_461  ))
// Xd_0__inst_mult_15_477  = CARRY(( (din_a[187] & din_b[182]) ) + ( Xd_0__inst_mult_15_462  ) + ( Xd_0__inst_mult_15_461  ))
// Xd_0__inst_mult_15_478  = SHARE((din_a[189] & din_b[181]))

	.dataa(!din_a[187]),
	.datab(!din_b[182]),
	.datac(!din_a[189]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_461 ),
	.sharein(Xd_0__inst_mult_15_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_476 ),
	.cout(Xd_0__inst_mult_15_477 ),
	.shareout(Xd_0__inst_mult_15_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_145 (
// Equation(s):
// Xd_0__inst_mult_15_480  = SUM(( (!din_a[186] & (((din_a[185] & din_b[184])))) # (din_a[186] & (!din_b[183] $ (((!din_a[185]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_466  ) + ( Xd_0__inst_mult_15_465  ))
// Xd_0__inst_mult_15_481  = CARRY(( (!din_a[186] & (((din_a[185] & din_b[184])))) # (din_a[186] & (!din_b[183] $ (((!din_a[185]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_466  ) + ( Xd_0__inst_mult_15_465  ))
// Xd_0__inst_mult_15_482  = SHARE((din_a[186] & (din_b[183] & (din_a[185] & din_b[184]))))

	.dataa(!din_a[186]),
	.datab(!din_b[183]),
	.datac(!din_a[185]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_465 ),
	.sharein(Xd_0__inst_mult_15_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_480 ),
	.cout(Xd_0__inst_mult_15_481 ),
	.shareout(Xd_0__inst_mult_15_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_67 (
// Equation(s):
// Xd_0__inst_mult_15_67_sumout  = SUM(( (din_a[189] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_68  = CARRY(( (din_a[189] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_69  = SHARE(GND)

	.dataa(!din_a[189]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_15_67_sumout ),
	.cout(Xd_0__inst_mult_15_68 ),
	.shareout(Xd_0__inst_mult_15_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_146 (
// Equation(s):
// Xd_0__inst_mult_15_484  = SUM(( (!din_a[183] & (((din_a[184] & din_b[185])))) # (din_a[183] & (!din_b[186] $ (((!din_a[184]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_15_470  ) + ( Xd_0__inst_mult_15_469  ))
// Xd_0__inst_mult_15_485  = CARRY(( (!din_a[183] & (((din_a[184] & din_b[185])))) # (din_a[183] & (!din_b[186] $ (((!din_a[184]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_15_470  ) + ( Xd_0__inst_mult_15_469  ))
// Xd_0__inst_mult_15_486  = SHARE((din_a[183] & (din_b[186] & (din_a[184] & din_b[185]))))

	.dataa(!din_a[183]),
	.datab(!din_b[186]),
	.datac(!din_a[184]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_469 ),
	.sharein(Xd_0__inst_mult_15_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_484 ),
	.cout(Xd_0__inst_mult_15_485 ),
	.shareout(Xd_0__inst_mult_15_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_147 (
// Equation(s):
// Xd_0__inst_mult_15_488  = SUM(( (din_a[180] & din_b[189]) ) + ( Xd_0__inst_mult_15_578  ) + ( Xd_0__inst_mult_15_577  ))
// Xd_0__inst_mult_15_489  = CARRY(( (din_a[180] & din_b[189]) ) + ( Xd_0__inst_mult_15_578  ) + ( Xd_0__inst_mult_15_577  ))
// Xd_0__inst_mult_15_490  = SHARE((din_a[180] & din_b[190]))

	.dataa(!din_a[180]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_577 ),
	.sharein(Xd_0__inst_mult_15_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_488 ),
	.cout(Xd_0__inst_mult_15_489 ),
	.shareout(Xd_0__inst_mult_15_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_133 (
// Equation(s):
// Xd_0__inst_mult_10_444  = SUM(( (din_a[127] & din_b[122]) ) + ( Xd_0__inst_mult_10_430  ) + ( Xd_0__inst_mult_10_429  ))
// Xd_0__inst_mult_10_445  = CARRY(( (din_a[127] & din_b[122]) ) + ( Xd_0__inst_mult_10_430  ) + ( Xd_0__inst_mult_10_429  ))
// Xd_0__inst_mult_10_446  = SHARE((din_a[129] & din_b[121]))

	.dataa(!din_a[127]),
	.datab(!din_b[122]),
	.datac(!din_a[129]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_429 ),
	.sharein(Xd_0__inst_mult_10_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_444 ),
	.cout(Xd_0__inst_mult_10_445 ),
	.shareout(Xd_0__inst_mult_10_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_134 (
// Equation(s):
// Xd_0__inst_mult_10_448  = SUM(( (!din_a[126] & (((din_a[125] & din_b[124])))) # (din_a[126] & (!din_b[123] $ (((!din_a[125]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_434  ) + ( Xd_0__inst_mult_10_433  ))
// Xd_0__inst_mult_10_449  = CARRY(( (!din_a[126] & (((din_a[125] & din_b[124])))) # (din_a[126] & (!din_b[123] $ (((!din_a[125]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_434  ) + ( Xd_0__inst_mult_10_433  ))
// Xd_0__inst_mult_10_450  = SHARE((din_a[126] & (din_b[123] & (din_a[125] & din_b[124]))))

	.dataa(!din_a[126]),
	.datab(!din_b[123]),
	.datac(!din_a[125]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_433 ),
	.sharein(Xd_0__inst_mult_10_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_448 ),
	.cout(Xd_0__inst_mult_10_449 ),
	.shareout(Xd_0__inst_mult_10_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_63 (
// Equation(s):
// Xd_0__inst_mult_10_63_sumout  = SUM(( (din_a[129] & din_b[120]) ) + ( Xd_0__inst_mult_11_69  ) + ( Xd_0__inst_mult_11_68  ))
// Xd_0__inst_mult_10_64  = CARRY(( (din_a[129] & din_b[120]) ) + ( Xd_0__inst_mult_11_69  ) + ( Xd_0__inst_mult_11_68  ))
// Xd_0__inst_mult_10_65  = SHARE(GND)

	.dataa(!din_a[129]),
	.datab(!din_b[120]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_68 ),
	.sharein(Xd_0__inst_mult_11_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_63_sumout ),
	.cout(Xd_0__inst_mult_10_64 ),
	.shareout(Xd_0__inst_mult_10_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_135 (
// Equation(s):
// Xd_0__inst_mult_10_452  = SUM(( (!din_a[123] & (((din_a[124] & din_b[125])))) # (din_a[123] & (!din_b[126] $ (((!din_a[124]) # (!din_b[125]))))) ) + ( Xd_0__inst_mult_10_438  ) + ( Xd_0__inst_mult_10_437  ))
// Xd_0__inst_mult_10_453  = CARRY(( (!din_a[123] & (((din_a[124] & din_b[125])))) # (din_a[123] & (!din_b[126] $ (((!din_a[124]) # (!din_b[125]))))) ) + ( Xd_0__inst_mult_10_438  ) + ( Xd_0__inst_mult_10_437  ))
// Xd_0__inst_mult_10_454  = SHARE((din_a[123] & (din_b[126] & (din_a[124] & din_b[125]))))

	.dataa(!din_a[123]),
	.datab(!din_b[126]),
	.datac(!din_a[124]),
	.datad(!din_b[125]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_437 ),
	.sharein(Xd_0__inst_mult_10_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_452 ),
	.cout(Xd_0__inst_mult_10_453 ),
	.shareout(Xd_0__inst_mult_10_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_136 (
// Equation(s):
// Xd_0__inst_mult_10_456  = SUM(( (din_a[120] & din_b[129]) ) + ( Xd_0__inst_mult_10_578  ) + ( Xd_0__inst_mult_10_577  ))
// Xd_0__inst_mult_10_457  = CARRY(( (din_a[120] & din_b[129]) ) + ( Xd_0__inst_mult_10_578  ) + ( Xd_0__inst_mult_10_577  ))
// Xd_0__inst_mult_10_458  = SHARE((din_a[120] & din_b[130]))

	.dataa(!din_a[120]),
	.datab(!din_b[129]),
	.datac(!din_b[130]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_577 ),
	.sharein(Xd_0__inst_mult_10_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_456 ),
	.cout(Xd_0__inst_mult_10_457 ),
	.shareout(Xd_0__inst_mult_10_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_137 (
// Equation(s):
// Xd_0__inst_mult_11_448  = SUM(( (din_a[139] & din_b[134]) ) + ( Xd_0__inst_mult_11_434  ) + ( Xd_0__inst_mult_11_433  ))
// Xd_0__inst_mult_11_449  = CARRY(( (din_a[139] & din_b[134]) ) + ( Xd_0__inst_mult_11_434  ) + ( Xd_0__inst_mult_11_433  ))
// Xd_0__inst_mult_11_450  = SHARE((din_a[141] & din_b[133]))

	.dataa(!din_a[139]),
	.datab(!din_b[134]),
	.datac(!din_a[141]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_433 ),
	.sharein(Xd_0__inst_mult_11_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_448 ),
	.cout(Xd_0__inst_mult_11_449 ),
	.shareout(Xd_0__inst_mult_11_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_138 (
// Equation(s):
// Xd_0__inst_mult_11_452  = SUM(( (!din_a[138] & (((din_a[137] & din_b[136])))) # (din_a[138] & (!din_b[135] $ (((!din_a[137]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_438  ) + ( Xd_0__inst_mult_11_437  ))
// Xd_0__inst_mult_11_453  = CARRY(( (!din_a[138] & (((din_a[137] & din_b[136])))) # (din_a[138] & (!din_b[135] $ (((!din_a[137]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_438  ) + ( Xd_0__inst_mult_11_437  ))
// Xd_0__inst_mult_11_454  = SHARE((din_a[138] & (din_b[135] & (din_a[137] & din_b[136]))))

	.dataa(!din_a[138]),
	.datab(!din_b[135]),
	.datac(!din_a[137]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_437 ),
	.sharein(Xd_0__inst_mult_11_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_452 ),
	.cout(Xd_0__inst_mult_11_453 ),
	.shareout(Xd_0__inst_mult_11_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_67 (
// Equation(s):
// Xd_0__inst_mult_11_67_sumout  = SUM(( (din_a[141] & din_b[132]) ) + ( Xd_0__inst_mult_8_69  ) + ( Xd_0__inst_mult_8_68  ))
// Xd_0__inst_mult_11_68  = CARRY(( (din_a[141] & din_b[132]) ) + ( Xd_0__inst_mult_8_69  ) + ( Xd_0__inst_mult_8_68  ))
// Xd_0__inst_mult_11_69  = SHARE(GND)

	.dataa(!din_a[141]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_68 ),
	.sharein(Xd_0__inst_mult_8_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_67_sumout ),
	.cout(Xd_0__inst_mult_11_68 ),
	.shareout(Xd_0__inst_mult_11_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_139 (
// Equation(s):
// Xd_0__inst_mult_11_456  = SUM(( (!din_a[135] & (((din_a[136] & din_b[137])))) # (din_a[135] & (!din_b[138] $ (((!din_a[136]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_11_442  ) + ( Xd_0__inst_mult_11_441  ))
// Xd_0__inst_mult_11_457  = CARRY(( (!din_a[135] & (((din_a[136] & din_b[137])))) # (din_a[135] & (!din_b[138] $ (((!din_a[136]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_11_442  ) + ( Xd_0__inst_mult_11_441  ))
// Xd_0__inst_mult_11_458  = SHARE((din_a[135] & (din_b[138] & (din_a[136] & din_b[137]))))

	.dataa(!din_a[135]),
	.datab(!din_b[138]),
	.datac(!din_a[136]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_441 ),
	.sharein(Xd_0__inst_mult_11_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_456 ),
	.cout(Xd_0__inst_mult_11_457 ),
	.shareout(Xd_0__inst_mult_11_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_140 (
// Equation(s):
// Xd_0__inst_mult_11_460  = SUM(( (din_a[132] & din_b[141]) ) + ( Xd_0__inst_mult_11_582  ) + ( Xd_0__inst_mult_11_581  ))
// Xd_0__inst_mult_11_461  = CARRY(( (din_a[132] & din_b[141]) ) + ( Xd_0__inst_mult_11_582  ) + ( Xd_0__inst_mult_11_581  ))
// Xd_0__inst_mult_11_462  = SHARE((din_a[132] & din_b[142]))

	.dataa(!din_a[132]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_581 ),
	.sharein(Xd_0__inst_mult_11_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_460 ),
	.cout(Xd_0__inst_mult_11_461 ),
	.shareout(Xd_0__inst_mult_11_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_137 (
// Equation(s):
// Xd_0__inst_mult_8_448  = SUM(( (din_a[103] & din_b[98]) ) + ( Xd_0__inst_mult_8_434  ) + ( Xd_0__inst_mult_8_433  ))
// Xd_0__inst_mult_8_449  = CARRY(( (din_a[103] & din_b[98]) ) + ( Xd_0__inst_mult_8_434  ) + ( Xd_0__inst_mult_8_433  ))
// Xd_0__inst_mult_8_450  = SHARE((din_a[105] & din_b[97]))

	.dataa(!din_a[103]),
	.datab(!din_b[98]),
	.datac(!din_a[105]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_433 ),
	.sharein(Xd_0__inst_mult_8_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_448 ),
	.cout(Xd_0__inst_mult_8_449 ),
	.shareout(Xd_0__inst_mult_8_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_138 (
// Equation(s):
// Xd_0__inst_mult_8_452  = SUM(( (!din_a[102] & (((din_a[101] & din_b[100])))) # (din_a[102] & (!din_b[99] $ (((!din_a[101]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_438  ) + ( Xd_0__inst_mult_8_437  ))
// Xd_0__inst_mult_8_453  = CARRY(( (!din_a[102] & (((din_a[101] & din_b[100])))) # (din_a[102] & (!din_b[99] $ (((!din_a[101]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_438  ) + ( Xd_0__inst_mult_8_437  ))
// Xd_0__inst_mult_8_454  = SHARE((din_a[102] & (din_b[99] & (din_a[101] & din_b[100]))))

	.dataa(!din_a[102]),
	.datab(!din_b[99]),
	.datac(!din_a[101]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_437 ),
	.sharein(Xd_0__inst_mult_8_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_452 ),
	.cout(Xd_0__inst_mult_8_453 ),
	.shareout(Xd_0__inst_mult_8_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_67 (
// Equation(s):
// Xd_0__inst_mult_8_67_sumout  = SUM(( (din_a[105] & din_b[96]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_68  = CARRY(( (din_a[105] & din_b[96]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_69  = SHARE(GND)

	.dataa(!din_a[105]),
	.datab(!din_b[96]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_8_67_sumout ),
	.cout(Xd_0__inst_mult_8_68 ),
	.shareout(Xd_0__inst_mult_8_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_139 (
// Equation(s):
// Xd_0__inst_mult_8_456  = SUM(( (!din_a[99] & (((din_a[100] & din_b[101])))) # (din_a[99] & (!din_b[102] $ (((!din_a[100]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_8_442  ) + ( Xd_0__inst_mult_8_441  ))
// Xd_0__inst_mult_8_457  = CARRY(( (!din_a[99] & (((din_a[100] & din_b[101])))) # (din_a[99] & (!din_b[102] $ (((!din_a[100]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_8_442  ) + ( Xd_0__inst_mult_8_441  ))
// Xd_0__inst_mult_8_458  = SHARE((din_a[99] & (din_b[102] & (din_a[100] & din_b[101]))))

	.dataa(!din_a[99]),
	.datab(!din_b[102]),
	.datac(!din_a[100]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_441 ),
	.sharein(Xd_0__inst_mult_8_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_456 ),
	.cout(Xd_0__inst_mult_8_457 ),
	.shareout(Xd_0__inst_mult_8_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_140 (
// Equation(s):
// Xd_0__inst_mult_8_460  = SUM(( (din_a[96] & din_b[105]) ) + ( Xd_0__inst_mult_8_582  ) + ( Xd_0__inst_mult_8_581  ))
// Xd_0__inst_mult_8_461  = CARRY(( (din_a[96] & din_b[105]) ) + ( Xd_0__inst_mult_8_582  ) + ( Xd_0__inst_mult_8_581  ))
// Xd_0__inst_mult_8_462  = SHARE((din_a[96] & din_b[106]))

	.dataa(!din_a[96]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_581 ),
	.sharein(Xd_0__inst_mult_8_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_460 ),
	.cout(Xd_0__inst_mult_8_461 ),
	.shareout(Xd_0__inst_mult_8_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_133 (
// Equation(s):
// Xd_0__inst_mult_9_444  = SUM(( (din_a[115] & din_b[110]) ) + ( Xd_0__inst_mult_9_430  ) + ( Xd_0__inst_mult_9_429  ))
// Xd_0__inst_mult_9_445  = CARRY(( (din_a[115] & din_b[110]) ) + ( Xd_0__inst_mult_9_430  ) + ( Xd_0__inst_mult_9_429  ))
// Xd_0__inst_mult_9_446  = SHARE((din_a[117] & din_b[109]))

	.dataa(!din_a[115]),
	.datab(!din_b[110]),
	.datac(!din_a[117]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_429 ),
	.sharein(Xd_0__inst_mult_9_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_444 ),
	.cout(Xd_0__inst_mult_9_445 ),
	.shareout(Xd_0__inst_mult_9_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_134 (
// Equation(s):
// Xd_0__inst_mult_9_448  = SUM(( (!din_a[114] & (((din_a[113] & din_b[112])))) # (din_a[114] & (!din_b[111] $ (((!din_a[113]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_434  ) + ( Xd_0__inst_mult_9_433  ))
// Xd_0__inst_mult_9_449  = CARRY(( (!din_a[114] & (((din_a[113] & din_b[112])))) # (din_a[114] & (!din_b[111] $ (((!din_a[113]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_434  ) + ( Xd_0__inst_mult_9_433  ))
// Xd_0__inst_mult_9_450  = SHARE((din_a[114] & (din_b[111] & (din_a[113] & din_b[112]))))

	.dataa(!din_a[114]),
	.datab(!din_b[111]),
	.datac(!din_a[113]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_433 ),
	.sharein(Xd_0__inst_mult_9_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_448 ),
	.cout(Xd_0__inst_mult_9_449 ),
	.shareout(Xd_0__inst_mult_9_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_135 (
// Equation(s):
// Xd_0__inst_mult_9_452  = SUM(( (!din_a[111] & (((din_a[112] & din_b[113])))) # (din_a[111] & (!din_b[114] $ (((!din_a[112]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_9_438  ) + ( Xd_0__inst_mult_9_437  ))
// Xd_0__inst_mult_9_453  = CARRY(( (!din_a[111] & (((din_a[112] & din_b[113])))) # (din_a[111] & (!din_b[114] $ (((!din_a[112]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_9_438  ) + ( Xd_0__inst_mult_9_437  ))
// Xd_0__inst_mult_9_454  = SHARE((din_a[111] & (din_b[114] & (din_a[112] & din_b[113]))))

	.dataa(!din_a[111]),
	.datab(!din_b[114]),
	.datac(!din_a[112]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_437 ),
	.sharein(Xd_0__inst_mult_9_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_452 ),
	.cout(Xd_0__inst_mult_9_453 ),
	.shareout(Xd_0__inst_mult_9_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_136 (
// Equation(s):
// Xd_0__inst_mult_9_456  = SUM(( (din_a[108] & din_b[117]) ) + ( Xd_0__inst_mult_9_578  ) + ( Xd_0__inst_mult_9_577  ))
// Xd_0__inst_mult_9_457  = CARRY(( (din_a[108] & din_b[117]) ) + ( Xd_0__inst_mult_9_578  ) + ( Xd_0__inst_mult_9_577  ))
// Xd_0__inst_mult_9_458  = SHARE((din_a[108] & din_b[118]))

	.dataa(!din_a[108]),
	.datab(!din_b[117]),
	.datac(!din_b[118]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_577 ),
	.sharein(Xd_0__inst_mult_9_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_456 ),
	.cout(Xd_0__inst_mult_9_457 ),
	.shareout(Xd_0__inst_mult_9_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_133 (
// Equation(s):
// Xd_0__inst_mult_6_444  = SUM(( (din_a[79] & din_b[74]) ) + ( Xd_0__inst_mult_6_430  ) + ( Xd_0__inst_mult_6_429  ))
// Xd_0__inst_mult_6_445  = CARRY(( (din_a[79] & din_b[74]) ) + ( Xd_0__inst_mult_6_430  ) + ( Xd_0__inst_mult_6_429  ))
// Xd_0__inst_mult_6_446  = SHARE((din_a[81] & din_b[73]))

	.dataa(!din_a[79]),
	.datab(!din_b[74]),
	.datac(!din_a[81]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_429 ),
	.sharein(Xd_0__inst_mult_6_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_444 ),
	.cout(Xd_0__inst_mult_6_445 ),
	.shareout(Xd_0__inst_mult_6_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_134 (
// Equation(s):
// Xd_0__inst_mult_6_448  = SUM(( (!din_a[78] & (((din_a[77] & din_b[76])))) # (din_a[78] & (!din_b[75] $ (((!din_a[77]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_434  ) + ( Xd_0__inst_mult_6_433  ))
// Xd_0__inst_mult_6_449  = CARRY(( (!din_a[78] & (((din_a[77] & din_b[76])))) # (din_a[78] & (!din_b[75] $ (((!din_a[77]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_434  ) + ( Xd_0__inst_mult_6_433  ))
// Xd_0__inst_mult_6_450  = SHARE((din_a[78] & (din_b[75] & (din_a[77] & din_b[76]))))

	.dataa(!din_a[78]),
	.datab(!din_b[75]),
	.datac(!din_a[77]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_433 ),
	.sharein(Xd_0__inst_mult_6_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_448 ),
	.cout(Xd_0__inst_mult_6_449 ),
	.shareout(Xd_0__inst_mult_6_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_63 (
// Equation(s):
// Xd_0__inst_mult_6_63_sumout  = SUM(( (din_a[81] & din_b[72]) ) + ( Xd_0__inst_mult_7_65  ) + ( Xd_0__inst_mult_7_64  ))
// Xd_0__inst_mult_6_64  = CARRY(( (din_a[81] & din_b[72]) ) + ( Xd_0__inst_mult_7_65  ) + ( Xd_0__inst_mult_7_64  ))
// Xd_0__inst_mult_6_65  = SHARE(GND)

	.dataa(!din_a[81]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_64 ),
	.sharein(Xd_0__inst_mult_7_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_63_sumout ),
	.cout(Xd_0__inst_mult_6_64 ),
	.shareout(Xd_0__inst_mult_6_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_135 (
// Equation(s):
// Xd_0__inst_mult_6_452  = SUM(( (!din_a[75] & (((din_a[76] & din_b[77])))) # (din_a[75] & (!din_b[78] $ (((!din_a[76]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_438  ) + ( Xd_0__inst_mult_6_437  ))
// Xd_0__inst_mult_6_453  = CARRY(( (!din_a[75] & (((din_a[76] & din_b[77])))) # (din_a[75] & (!din_b[78] $ (((!din_a[76]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_438  ) + ( Xd_0__inst_mult_6_437  ))
// Xd_0__inst_mult_6_454  = SHARE((din_a[75] & (din_b[78] & (din_a[76] & din_b[77]))))

	.dataa(!din_a[75]),
	.datab(!din_b[78]),
	.datac(!din_a[76]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_437 ),
	.sharein(Xd_0__inst_mult_6_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_452 ),
	.cout(Xd_0__inst_mult_6_453 ),
	.shareout(Xd_0__inst_mult_6_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_136 (
// Equation(s):
// Xd_0__inst_mult_6_456  = SUM(( (din_a[72] & din_b[81]) ) + ( Xd_0__inst_mult_6_578  ) + ( Xd_0__inst_mult_6_577  ))
// Xd_0__inst_mult_6_457  = CARRY(( (din_a[72] & din_b[81]) ) + ( Xd_0__inst_mult_6_578  ) + ( Xd_0__inst_mult_6_577  ))
// Xd_0__inst_mult_6_458  = SHARE((din_a[72] & din_b[82]))

	.dataa(!din_a[72]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_577 ),
	.sharein(Xd_0__inst_mult_6_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_456 ),
	.cout(Xd_0__inst_mult_6_457 ),
	.shareout(Xd_0__inst_mult_6_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_129 (
// Equation(s):
// Xd_0__inst_mult_7_428  = SUM(( (din_a[91] & din_b[86]) ) + ( Xd_0__inst_mult_7_414  ) + ( Xd_0__inst_mult_7_413  ))
// Xd_0__inst_mult_7_429  = CARRY(( (din_a[91] & din_b[86]) ) + ( Xd_0__inst_mult_7_414  ) + ( Xd_0__inst_mult_7_413  ))
// Xd_0__inst_mult_7_430  = SHARE((din_a[93] & din_b[85]))

	.dataa(!din_a[91]),
	.datab(!din_b[86]),
	.datac(!din_a[93]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_413 ),
	.sharein(Xd_0__inst_mult_7_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_428 ),
	.cout(Xd_0__inst_mult_7_429 ),
	.shareout(Xd_0__inst_mult_7_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_130 (
// Equation(s):
// Xd_0__inst_mult_7_432  = SUM(( (!din_a[90] & (((din_a[89] & din_b[88])))) # (din_a[90] & (!din_b[87] $ (((!din_a[89]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_418  ) + ( Xd_0__inst_mult_7_417  ))
// Xd_0__inst_mult_7_433  = CARRY(( (!din_a[90] & (((din_a[89] & din_b[88])))) # (din_a[90] & (!din_b[87] $ (((!din_a[89]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_418  ) + ( Xd_0__inst_mult_7_417  ))
// Xd_0__inst_mult_7_434  = SHARE((din_a[90] & (din_b[87] & (din_a[89] & din_b[88]))))

	.dataa(!din_a[90]),
	.datab(!din_b[87]),
	.datac(!din_a[89]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_417 ),
	.sharein(Xd_0__inst_mult_7_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_432 ),
	.cout(Xd_0__inst_mult_7_433 ),
	.shareout(Xd_0__inst_mult_7_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_63 (
// Equation(s):
// Xd_0__inst_mult_7_63_sumout  = SUM(( (din_a[93] & din_b[84]) ) + ( Xd_0__inst_mult_4_69  ) + ( Xd_0__inst_mult_4_68  ))
// Xd_0__inst_mult_7_64  = CARRY(( (din_a[93] & din_b[84]) ) + ( Xd_0__inst_mult_4_69  ) + ( Xd_0__inst_mult_4_68  ))
// Xd_0__inst_mult_7_65  = SHARE(GND)

	.dataa(!din_a[93]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_68 ),
	.sharein(Xd_0__inst_mult_4_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_63_sumout ),
	.cout(Xd_0__inst_mult_7_64 ),
	.shareout(Xd_0__inst_mult_7_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_131 (
// Equation(s):
// Xd_0__inst_mult_7_436  = SUM(( (!din_a[87] & (((din_a[88] & din_b[89])))) # (din_a[87] & (!din_b[90] $ (((!din_a[88]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_422  ) + ( Xd_0__inst_mult_7_421  ))
// Xd_0__inst_mult_7_437  = CARRY(( (!din_a[87] & (((din_a[88] & din_b[89])))) # (din_a[87] & (!din_b[90] $ (((!din_a[88]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_422  ) + ( Xd_0__inst_mult_7_421  ))
// Xd_0__inst_mult_7_438  = SHARE((din_a[87] & (din_b[90] & (din_a[88] & din_b[89]))))

	.dataa(!din_a[87]),
	.datab(!din_b[90]),
	.datac(!din_a[88]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_421 ),
	.sharein(Xd_0__inst_mult_7_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_436 ),
	.cout(Xd_0__inst_mult_7_437 ),
	.shareout(Xd_0__inst_mult_7_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_132 (
// Equation(s):
// Xd_0__inst_mult_7_440  = SUM(( (din_a[84] & din_b[93]) ) + ( Xd_0__inst_mult_7_578  ) + ( Xd_0__inst_mult_7_577  ))
// Xd_0__inst_mult_7_441  = CARRY(( (din_a[84] & din_b[93]) ) + ( Xd_0__inst_mult_7_578  ) + ( Xd_0__inst_mult_7_577  ))
// Xd_0__inst_mult_7_442  = SHARE((din_a[84] & din_b[94]))

	.dataa(!din_a[84]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_577 ),
	.sharein(Xd_0__inst_mult_7_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_440 ),
	.cout(Xd_0__inst_mult_7_441 ),
	.shareout(Xd_0__inst_mult_7_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_142 (
// Equation(s):
// Xd_0__inst_mult_4_468  = SUM(( (din_a[55] & din_b[50]) ) + ( Xd_0__inst_mult_4_454  ) + ( Xd_0__inst_mult_4_453  ))
// Xd_0__inst_mult_4_469  = CARRY(( (din_a[55] & din_b[50]) ) + ( Xd_0__inst_mult_4_454  ) + ( Xd_0__inst_mult_4_453  ))
// Xd_0__inst_mult_4_470  = SHARE((din_a[57] & din_b[49]))

	.dataa(!din_a[55]),
	.datab(!din_b[50]),
	.datac(!din_a[57]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_453 ),
	.sharein(Xd_0__inst_mult_4_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_468 ),
	.cout(Xd_0__inst_mult_4_469 ),
	.shareout(Xd_0__inst_mult_4_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_143 (
// Equation(s):
// Xd_0__inst_mult_4_472  = SUM(( (!din_a[54] & (((din_a[53] & din_b[52])))) # (din_a[54] & (!din_b[51] $ (((!din_a[53]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_458  ) + ( Xd_0__inst_mult_4_457  ))
// Xd_0__inst_mult_4_473  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[52])))) # (din_a[54] & (!din_b[51] $ (((!din_a[53]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_458  ) + ( Xd_0__inst_mult_4_457  ))
// Xd_0__inst_mult_4_474  = SHARE((din_a[54] & (din_b[51] & (din_a[53] & din_b[52]))))

	.dataa(!din_a[54]),
	.datab(!din_b[51]),
	.datac(!din_a[53]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_457 ),
	.sharein(Xd_0__inst_mult_4_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_472 ),
	.cout(Xd_0__inst_mult_4_473 ),
	.shareout(Xd_0__inst_mult_4_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_67 (
// Equation(s):
// Xd_0__inst_mult_4_67_sumout  = SUM(( (din_a[57] & din_b[48]) ) + ( Xd_0__inst_mult_3_49  ) + ( Xd_0__inst_mult_3_48  ))
// Xd_0__inst_mult_4_68  = CARRY(( (din_a[57] & din_b[48]) ) + ( Xd_0__inst_mult_3_49  ) + ( Xd_0__inst_mult_3_48  ))
// Xd_0__inst_mult_4_69  = SHARE(GND)

	.dataa(!din_a[57]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_48 ),
	.sharein(Xd_0__inst_mult_3_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_67_sumout ),
	.cout(Xd_0__inst_mult_4_68 ),
	.shareout(Xd_0__inst_mult_4_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_144 (
// Equation(s):
// Xd_0__inst_mult_4_476  = SUM(( (!din_a[51] & (((din_a[52] & din_b[53])))) # (din_a[51] & (!din_b[54] $ (((!din_a[52]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_462  ) + ( Xd_0__inst_mult_4_461  ))
// Xd_0__inst_mult_4_477  = CARRY(( (!din_a[51] & (((din_a[52] & din_b[53])))) # (din_a[51] & (!din_b[54] $ (((!din_a[52]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_462  ) + ( Xd_0__inst_mult_4_461  ))
// Xd_0__inst_mult_4_478  = SHARE((din_a[51] & (din_b[54] & (din_a[52] & din_b[53]))))

	.dataa(!din_a[51]),
	.datab(!din_b[54]),
	.datac(!din_a[52]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_461 ),
	.sharein(Xd_0__inst_mult_4_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_476 ),
	.cout(Xd_0__inst_mult_4_477 ),
	.shareout(Xd_0__inst_mult_4_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_145 (
// Equation(s):
// Xd_0__inst_mult_4_480  = SUM(( (din_a[48] & din_b[57]) ) + ( Xd_0__inst_mult_4_578  ) + ( Xd_0__inst_mult_4_577  ))
// Xd_0__inst_mult_4_481  = CARRY(( (din_a[48] & din_b[57]) ) + ( Xd_0__inst_mult_4_578  ) + ( Xd_0__inst_mult_4_577  ))
// Xd_0__inst_mult_4_482  = SHARE((din_a[48] & din_b[58]))

	.dataa(!din_a[48]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_577 ),
	.sharein(Xd_0__inst_mult_4_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_480 ),
	.cout(Xd_0__inst_mult_4_481 ),
	.shareout(Xd_0__inst_mult_4_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_129 (
// Equation(s):
// Xd_0__inst_mult_5_428  = SUM(( (din_a[67] & din_b[62]) ) + ( Xd_0__inst_mult_5_414  ) + ( Xd_0__inst_mult_5_413  ))
// Xd_0__inst_mult_5_429  = CARRY(( (din_a[67] & din_b[62]) ) + ( Xd_0__inst_mult_5_414  ) + ( Xd_0__inst_mult_5_413  ))
// Xd_0__inst_mult_5_430  = SHARE((din_a[69] & din_b[61]))

	.dataa(!din_a[67]),
	.datab(!din_b[62]),
	.datac(!din_a[69]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_413 ),
	.sharein(Xd_0__inst_mult_5_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_428 ),
	.cout(Xd_0__inst_mult_5_429 ),
	.shareout(Xd_0__inst_mult_5_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_130 (
// Equation(s):
// Xd_0__inst_mult_5_432  = SUM(( (!din_a[66] & (((din_a[65] & din_b[64])))) # (din_a[66] & (!din_b[63] $ (((!din_a[65]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_418  ) + ( Xd_0__inst_mult_5_417  ))
// Xd_0__inst_mult_5_433  = CARRY(( (!din_a[66] & (((din_a[65] & din_b[64])))) # (din_a[66] & (!din_b[63] $ (((!din_a[65]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_418  ) + ( Xd_0__inst_mult_5_417  ))
// Xd_0__inst_mult_5_434  = SHARE((din_a[66] & (din_b[63] & (din_a[65] & din_b[64]))))

	.dataa(!din_a[66]),
	.datab(!din_b[63]),
	.datac(!din_a[65]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_417 ),
	.sharein(Xd_0__inst_mult_5_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_432 ),
	.cout(Xd_0__inst_mult_5_433 ),
	.shareout(Xd_0__inst_mult_5_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_131 (
// Equation(s):
// Xd_0__inst_mult_5_436  = SUM(( (!din_a[63] & (((din_a[64] & din_b[65])))) # (din_a[63] & (!din_b[66] $ (((!din_a[64]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_422  ) + ( Xd_0__inst_mult_5_421  ))
// Xd_0__inst_mult_5_437  = CARRY(( (!din_a[63] & (((din_a[64] & din_b[65])))) # (din_a[63] & (!din_b[66] $ (((!din_a[64]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_422  ) + ( Xd_0__inst_mult_5_421  ))
// Xd_0__inst_mult_5_438  = SHARE((din_a[63] & (din_b[66] & (din_a[64] & din_b[65]))))

	.dataa(!din_a[63]),
	.datab(!din_b[66]),
	.datac(!din_a[64]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_421 ),
	.sharein(Xd_0__inst_mult_5_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_436 ),
	.cout(Xd_0__inst_mult_5_437 ),
	.shareout(Xd_0__inst_mult_5_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_132 (
// Equation(s):
// Xd_0__inst_mult_5_440  = SUM(( (din_a[60] & din_b[69]) ) + ( Xd_0__inst_mult_5_578  ) + ( Xd_0__inst_mult_5_577  ))
// Xd_0__inst_mult_5_441  = CARRY(( (din_a[60] & din_b[69]) ) + ( Xd_0__inst_mult_5_578  ) + ( Xd_0__inst_mult_5_577  ))
// Xd_0__inst_mult_5_442  = SHARE((din_a[60] & din_b[70]))

	.dataa(!din_a[60]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_577 ),
	.sharein(Xd_0__inst_mult_5_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_440 ),
	.cout(Xd_0__inst_mult_5_441 ),
	.shareout(Xd_0__inst_mult_5_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_133 (
// Equation(s):
// Xd_0__inst_mult_2_432  = SUM(( (din_a[31] & din_b[26]) ) + ( Xd_0__inst_mult_2_418  ) + ( Xd_0__inst_mult_2_417  ))
// Xd_0__inst_mult_2_433  = CARRY(( (din_a[31] & din_b[26]) ) + ( Xd_0__inst_mult_2_418  ) + ( Xd_0__inst_mult_2_417  ))
// Xd_0__inst_mult_2_434  = SHARE((din_a[33] & din_b[25]))

	.dataa(!din_a[31]),
	.datab(!din_b[26]),
	.datac(!din_a[33]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_417 ),
	.sharein(Xd_0__inst_mult_2_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_432 ),
	.cout(Xd_0__inst_mult_2_433 ),
	.shareout(Xd_0__inst_mult_2_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_134 (
// Equation(s):
// Xd_0__inst_mult_2_436  = SUM(( (!din_a[30] & (((din_a[29] & din_b[28])))) # (din_a[30] & (!din_b[27] $ (((!din_a[29]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_422  ) + ( Xd_0__inst_mult_2_421  ))
// Xd_0__inst_mult_2_437  = CARRY(( (!din_a[30] & (((din_a[29] & din_b[28])))) # (din_a[30] & (!din_b[27] $ (((!din_a[29]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_422  ) + ( Xd_0__inst_mult_2_421  ))
// Xd_0__inst_mult_2_438  = SHARE((din_a[30] & (din_b[27] & (din_a[29] & din_b[28]))))

	.dataa(!din_a[30]),
	.datab(!din_b[27]),
	.datac(!din_a[29]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_421 ),
	.sharein(Xd_0__inst_mult_2_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_436 ),
	.cout(Xd_0__inst_mult_2_437 ),
	.shareout(Xd_0__inst_mult_2_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_135 (
// Equation(s):
// Xd_0__inst_mult_2_440  = SUM(( (!din_a[27] & (((din_a[28] & din_b[29])))) # (din_a[27] & (!din_b[30] $ (((!din_a[28]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_426  ) + ( Xd_0__inst_mult_2_425  ))
// Xd_0__inst_mult_2_441  = CARRY(( (!din_a[27] & (((din_a[28] & din_b[29])))) # (din_a[27] & (!din_b[30] $ (((!din_a[28]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_426  ) + ( Xd_0__inst_mult_2_425  ))
// Xd_0__inst_mult_2_442  = SHARE((din_a[27] & (din_b[30] & (din_a[28] & din_b[29]))))

	.dataa(!din_a[27]),
	.datab(!din_b[30]),
	.datac(!din_a[28]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_425 ),
	.sharein(Xd_0__inst_mult_2_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_440 ),
	.cout(Xd_0__inst_mult_2_441 ),
	.shareout(Xd_0__inst_mult_2_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_136 (
// Equation(s):
// Xd_0__inst_mult_2_444  = SUM(( (din_a[24] & din_b[33]) ) + ( Xd_0__inst_mult_2_582  ) + ( Xd_0__inst_mult_2_581  ))
// Xd_0__inst_mult_2_445  = CARRY(( (din_a[24] & din_b[33]) ) + ( Xd_0__inst_mult_2_582  ) + ( Xd_0__inst_mult_2_581  ))
// Xd_0__inst_mult_2_446  = SHARE((din_a[24] & din_b[34]))

	.dataa(!din_a[24]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_581 ),
	.sharein(Xd_0__inst_mult_2_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_444 ),
	.cout(Xd_0__inst_mult_2_445 ),
	.shareout(Xd_0__inst_mult_2_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_129 (
// Equation(s):
// Xd_0__inst_mult_3_428  = SUM(( (din_a[43] & din_b[38]) ) + ( Xd_0__inst_mult_3_414  ) + ( Xd_0__inst_mult_3_413  ))
// Xd_0__inst_mult_3_429  = CARRY(( (din_a[43] & din_b[38]) ) + ( Xd_0__inst_mult_3_414  ) + ( Xd_0__inst_mult_3_413  ))
// Xd_0__inst_mult_3_430  = SHARE((din_a[45] & din_b[37]))

	.dataa(!din_a[43]),
	.datab(!din_b[38]),
	.datac(!din_a[45]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_413 ),
	.sharein(Xd_0__inst_mult_3_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_428 ),
	.cout(Xd_0__inst_mult_3_429 ),
	.shareout(Xd_0__inst_mult_3_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_130 (
// Equation(s):
// Xd_0__inst_mult_3_432  = SUM(( (!din_a[42] & (((din_a[41] & din_b[40])))) # (din_a[42] & (!din_b[39] $ (((!din_a[41]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_418  ) + ( Xd_0__inst_mult_3_417  ))
// Xd_0__inst_mult_3_433  = CARRY(( (!din_a[42] & (((din_a[41] & din_b[40])))) # (din_a[42] & (!din_b[39] $ (((!din_a[41]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_418  ) + ( Xd_0__inst_mult_3_417  ))
// Xd_0__inst_mult_3_434  = SHARE((din_a[42] & (din_b[39] & (din_a[41] & din_b[40]))))

	.dataa(!din_a[42]),
	.datab(!din_b[39]),
	.datac(!din_a[41]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_417 ),
	.sharein(Xd_0__inst_mult_3_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_432 ),
	.cout(Xd_0__inst_mult_3_433 ),
	.shareout(Xd_0__inst_mult_3_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_131 (
// Equation(s):
// Xd_0__inst_mult_3_436  = SUM(( (!din_a[39] & (((din_a[40] & din_b[41])))) # (din_a[39] & (!din_b[42] $ (((!din_a[40]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_422  ) + ( Xd_0__inst_mult_3_421  ))
// Xd_0__inst_mult_3_437  = CARRY(( (!din_a[39] & (((din_a[40] & din_b[41])))) # (din_a[39] & (!din_b[42] $ (((!din_a[40]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_422  ) + ( Xd_0__inst_mult_3_421  ))
// Xd_0__inst_mult_3_438  = SHARE((din_a[39] & (din_b[42] & (din_a[40] & din_b[41]))))

	.dataa(!din_a[39]),
	.datab(!din_b[42]),
	.datac(!din_a[40]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_421 ),
	.sharein(Xd_0__inst_mult_3_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_436 ),
	.cout(Xd_0__inst_mult_3_437 ),
	.shareout(Xd_0__inst_mult_3_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_132 (
// Equation(s):
// Xd_0__inst_mult_3_440  = SUM(( (din_a[36] & din_b[45]) ) + ( Xd_0__inst_mult_3_578  ) + ( Xd_0__inst_mult_3_577  ))
// Xd_0__inst_mult_3_441  = CARRY(( (din_a[36] & din_b[45]) ) + ( Xd_0__inst_mult_3_578  ) + ( Xd_0__inst_mult_3_577  ))
// Xd_0__inst_mult_3_442  = SHARE((din_a[36] & din_b[46]))

	.dataa(!din_a[36]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_577 ),
	.sharein(Xd_0__inst_mult_3_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_440 ),
	.cout(Xd_0__inst_mult_3_441 ),
	.shareout(Xd_0__inst_mult_3_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_133 (
// Equation(s):
// Xd_0__inst_mult_0_432  = SUM(( (din_a[7] & din_b[2]) ) + ( Xd_0__inst_mult_0_418  ) + ( Xd_0__inst_mult_0_417  ))
// Xd_0__inst_mult_0_433  = CARRY(( (din_a[7] & din_b[2]) ) + ( Xd_0__inst_mult_0_418  ) + ( Xd_0__inst_mult_0_417  ))
// Xd_0__inst_mult_0_434  = SHARE((din_a[9] & din_b[1]))

	.dataa(!din_a[7]),
	.datab(!din_b[2]),
	.datac(!din_a[9]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_417 ),
	.sharein(Xd_0__inst_mult_0_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_432 ),
	.cout(Xd_0__inst_mult_0_433 ),
	.shareout(Xd_0__inst_mult_0_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_134 (
// Equation(s):
// Xd_0__inst_mult_0_436  = SUM(( (!din_a[6] & (((din_a[5] & din_b[4])))) # (din_a[6] & (!din_b[3] $ (((!din_a[5]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_422  ) + ( Xd_0__inst_mult_0_421  ))
// Xd_0__inst_mult_0_437  = CARRY(( (!din_a[6] & (((din_a[5] & din_b[4])))) # (din_a[6] & (!din_b[3] $ (((!din_a[5]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_422  ) + ( Xd_0__inst_mult_0_421  ))
// Xd_0__inst_mult_0_438  = SHARE((din_a[6] & (din_b[3] & (din_a[5] & din_b[4]))))

	.dataa(!din_a[6]),
	.datab(!din_b[3]),
	.datac(!din_a[5]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_421 ),
	.sharein(Xd_0__inst_mult_0_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_436 ),
	.cout(Xd_0__inst_mult_0_437 ),
	.shareout(Xd_0__inst_mult_0_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_135 (
// Equation(s):
// Xd_0__inst_mult_0_440  = SUM(( (!din_a[3] & (((din_a[4] & din_b[5])))) # (din_a[3] & (!din_b[6] $ (((!din_a[4]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_426  ) + ( Xd_0__inst_mult_0_425  ))
// Xd_0__inst_mult_0_441  = CARRY(( (!din_a[3] & (((din_a[4] & din_b[5])))) # (din_a[3] & (!din_b[6] $ (((!din_a[4]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_426  ) + ( Xd_0__inst_mult_0_425  ))
// Xd_0__inst_mult_0_442  = SHARE((din_a[3] & (din_b[6] & (din_a[4] & din_b[5]))))

	.dataa(!din_a[3]),
	.datab(!din_b[6]),
	.datac(!din_a[4]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_425 ),
	.sharein(Xd_0__inst_mult_0_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_440 ),
	.cout(Xd_0__inst_mult_0_441 ),
	.shareout(Xd_0__inst_mult_0_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_136 (
// Equation(s):
// Xd_0__inst_mult_0_444  = SUM(( (din_a[0] & din_b[9]) ) + ( Xd_0__inst_mult_0_582  ) + ( Xd_0__inst_mult_0_581  ))
// Xd_0__inst_mult_0_445  = CARRY(( (din_a[0] & din_b[9]) ) + ( Xd_0__inst_mult_0_582  ) + ( Xd_0__inst_mult_0_581  ))
// Xd_0__inst_mult_0_446  = SHARE((din_a[0] & din_b[10]))

	.dataa(!din_a[0]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_581 ),
	.sharein(Xd_0__inst_mult_0_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_444 ),
	.cout(Xd_0__inst_mult_0_445 ),
	.shareout(Xd_0__inst_mult_0_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_133 (
// Equation(s):
// Xd_0__inst_mult_1_432  = SUM(( (din_a[19] & din_b[14]) ) + ( Xd_0__inst_mult_1_418  ) + ( Xd_0__inst_mult_1_417  ))
// Xd_0__inst_mult_1_433  = CARRY(( (din_a[19] & din_b[14]) ) + ( Xd_0__inst_mult_1_418  ) + ( Xd_0__inst_mult_1_417  ))
// Xd_0__inst_mult_1_434  = SHARE((din_a[21] & din_b[13]))

	.dataa(!din_a[19]),
	.datab(!din_b[14]),
	.datac(!din_a[21]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_417 ),
	.sharein(Xd_0__inst_mult_1_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_432 ),
	.cout(Xd_0__inst_mult_1_433 ),
	.shareout(Xd_0__inst_mult_1_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_134 (
// Equation(s):
// Xd_0__inst_mult_1_436  = SUM(( (!din_a[18] & (((din_a[17] & din_b[16])))) # (din_a[18] & (!din_b[15] $ (((!din_a[17]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_422  ) + ( Xd_0__inst_mult_1_421  ))
// Xd_0__inst_mult_1_437  = CARRY(( (!din_a[18] & (((din_a[17] & din_b[16])))) # (din_a[18] & (!din_b[15] $ (((!din_a[17]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_422  ) + ( Xd_0__inst_mult_1_421  ))
// Xd_0__inst_mult_1_438  = SHARE((din_a[18] & (din_b[15] & (din_a[17] & din_b[16]))))

	.dataa(!din_a[18]),
	.datab(!din_b[15]),
	.datac(!din_a[17]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_421 ),
	.sharein(Xd_0__inst_mult_1_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_436 ),
	.cout(Xd_0__inst_mult_1_437 ),
	.shareout(Xd_0__inst_mult_1_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_135 (
// Equation(s):
// Xd_0__inst_mult_1_440  = SUM(( (!din_a[15] & (((din_a[16] & din_b[17])))) # (din_a[15] & (!din_b[18] $ (((!din_a[16]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_426  ) + ( Xd_0__inst_mult_1_425  ))
// Xd_0__inst_mult_1_441  = CARRY(( (!din_a[15] & (((din_a[16] & din_b[17])))) # (din_a[15] & (!din_b[18] $ (((!din_a[16]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_426  ) + ( Xd_0__inst_mult_1_425  ))
// Xd_0__inst_mult_1_442  = SHARE((din_a[15] & (din_b[18] & (din_a[16] & din_b[17]))))

	.dataa(!din_a[15]),
	.datab(!din_b[18]),
	.datac(!din_a[16]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_425 ),
	.sharein(Xd_0__inst_mult_1_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_440 ),
	.cout(Xd_0__inst_mult_1_441 ),
	.shareout(Xd_0__inst_mult_1_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_136 (
// Equation(s):
// Xd_0__inst_mult_1_444  = SUM(( (din_a[12] & din_b[21]) ) + ( Xd_0__inst_mult_1_582  ) + ( Xd_0__inst_mult_1_581  ))
// Xd_0__inst_mult_1_445  = CARRY(( (din_a[12] & din_b[21]) ) + ( Xd_0__inst_mult_1_582  ) + ( Xd_0__inst_mult_1_581  ))
// Xd_0__inst_mult_1_446  = SHARE((din_a[12] & din_b[22]))

	.dataa(!din_a[12]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_581 ),
	.sharein(Xd_0__inst_mult_1_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_444 ),
	.cout(Xd_0__inst_mult_1_445 ),
	.shareout(Xd_0__inst_mult_1_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_144 (
// Equation(s):
// Xd_0__inst_mult_12_488  = SUM(( (din_a[152] & din_b[146]) ) + ( Xd_0__inst_mult_12_474  ) + ( Xd_0__inst_mult_12_473  ))
// Xd_0__inst_mult_12_489  = CARRY(( (din_a[152] & din_b[146]) ) + ( Xd_0__inst_mult_12_474  ) + ( Xd_0__inst_mult_12_473  ))
// Xd_0__inst_mult_12_490  = SHARE((din_a[154] & din_b[145]))

	.dataa(!din_a[152]),
	.datab(!din_b[146]),
	.datac(!din_a[154]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_473 ),
	.sharein(Xd_0__inst_mult_12_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_488 ),
	.cout(Xd_0__inst_mult_12_489 ),
	.shareout(Xd_0__inst_mult_12_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_145 (
// Equation(s):
// Xd_0__inst_mult_12_492  = SUM(( (!din_a[151] & (((din_a[150] & din_b[148])))) # (din_a[151] & (!din_b[147] $ (((!din_a[150]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_478  ) + ( Xd_0__inst_mult_12_477  ))
// Xd_0__inst_mult_12_493  = CARRY(( (!din_a[151] & (((din_a[150] & din_b[148])))) # (din_a[151] & (!din_b[147] $ (((!din_a[150]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_478  ) + ( Xd_0__inst_mult_12_477  ))
// Xd_0__inst_mult_12_494  = SHARE((din_a[151] & (din_b[147] & (din_a[150] & din_b[148]))))

	.dataa(!din_a[151]),
	.datab(!din_b[147]),
	.datac(!din_a[150]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_477 ),
	.sharein(Xd_0__inst_mult_12_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_492 ),
	.cout(Xd_0__inst_mult_12_493 ),
	.shareout(Xd_0__inst_mult_12_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_146 (
// Equation(s):
// Xd_0__inst_mult_12_496  = SUM(( (din_a[149] & din_b[149]) ) + ( Xd_0__inst_mult_12_482  ) + ( Xd_0__inst_mult_12_481  ))
// Xd_0__inst_mult_12_497  = CARRY(( (din_a[149] & din_b[149]) ) + ( Xd_0__inst_mult_12_482  ) + ( Xd_0__inst_mult_12_481  ))
// Xd_0__inst_mult_12_498  = SHARE((din_a[149] & din_b[150]))

	.dataa(!din_a[149]),
	.datab(!din_b[149]),
	.datac(!din_b[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_481 ),
	.sharein(Xd_0__inst_mult_12_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_496 ),
	.cout(Xd_0__inst_mult_12_497 ),
	.shareout(Xd_0__inst_mult_12_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_147 (
// Equation(s):
// Xd_0__inst_mult_12_500  = SUM(( (din_a[145] & din_b[153]) ) + ( Xd_0__inst_mult_12_486  ) + ( Xd_0__inst_mult_12_485  ))
// Xd_0__inst_mult_12_501  = CARRY(( (din_a[145] & din_b[153]) ) + ( Xd_0__inst_mult_12_486  ) + ( Xd_0__inst_mult_12_485  ))
// Xd_0__inst_mult_12_502  = SHARE((din_a[145] & din_b[154]))

	.dataa(!din_a[145]),
	.datab(!din_b[153]),
	.datac(!din_b[154]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_485 ),
	.sharein(Xd_0__inst_mult_12_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_500 ),
	.cout(Xd_0__inst_mult_12_501 ),
	.shareout(Xd_0__inst_mult_12_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_148 (
// Equation(s):
// Xd_0__inst_mult_12_504  = SUM(( (!din_a[147] & (((din_a[146] & din_b[152])))) # (din_a[147] & (!din_b[151] $ (((!din_a[146]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_578  ) + ( Xd_0__inst_mult_12_577  ))
// Xd_0__inst_mult_12_505  = CARRY(( (!din_a[147] & (((din_a[146] & din_b[152])))) # (din_a[147] & (!din_b[151] $ (((!din_a[146]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_578  ) + ( Xd_0__inst_mult_12_577  ))
// Xd_0__inst_mult_12_506  = SHARE((din_a[147] & (din_b[151] & (din_a[146] & din_b[152]))))

	.dataa(!din_a[147]),
	.datab(!din_b[151]),
	.datac(!din_a[146]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_577 ),
	.sharein(Xd_0__inst_mult_12_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_504 ),
	.cout(Xd_0__inst_mult_12_505 ),
	.shareout(Xd_0__inst_mult_12_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_141 (
// Equation(s):
// Xd_0__inst_mult_13_464  = SUM(( (din_a[164] & din_b[158]) ) + ( Xd_0__inst_mult_13_450  ) + ( Xd_0__inst_mult_13_449  ))
// Xd_0__inst_mult_13_465  = CARRY(( (din_a[164] & din_b[158]) ) + ( Xd_0__inst_mult_13_450  ) + ( Xd_0__inst_mult_13_449  ))
// Xd_0__inst_mult_13_466  = SHARE((din_a[166] & din_b[157]))

	.dataa(!din_a[164]),
	.datab(!din_b[158]),
	.datac(!din_a[166]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_449 ),
	.sharein(Xd_0__inst_mult_13_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_464 ),
	.cout(Xd_0__inst_mult_13_465 ),
	.shareout(Xd_0__inst_mult_13_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_142 (
// Equation(s):
// Xd_0__inst_mult_13_468  = SUM(( (!din_a[163] & (((din_a[162] & din_b[160])))) # (din_a[163] & (!din_b[159] $ (((!din_a[162]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_454  ) + ( Xd_0__inst_mult_13_453  ))
// Xd_0__inst_mult_13_469  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[160])))) # (din_a[163] & (!din_b[159] $ (((!din_a[162]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_454  ) + ( Xd_0__inst_mult_13_453  ))
// Xd_0__inst_mult_13_470  = SHARE((din_a[163] & (din_b[159] & (din_a[162] & din_b[160]))))

	.dataa(!din_a[163]),
	.datab(!din_b[159]),
	.datac(!din_a[162]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_453 ),
	.sharein(Xd_0__inst_mult_13_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_468 ),
	.cout(Xd_0__inst_mult_13_469 ),
	.shareout(Xd_0__inst_mult_13_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_143 (
// Equation(s):
// Xd_0__inst_mult_13_472  = SUM(( (din_a[161] & din_b[161]) ) + ( Xd_0__inst_mult_13_458  ) + ( Xd_0__inst_mult_13_457  ))
// Xd_0__inst_mult_13_473  = CARRY(( (din_a[161] & din_b[161]) ) + ( Xd_0__inst_mult_13_458  ) + ( Xd_0__inst_mult_13_457  ))
// Xd_0__inst_mult_13_474  = SHARE((din_a[161] & din_b[162]))

	.dataa(!din_a[161]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_457 ),
	.sharein(Xd_0__inst_mult_13_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_472 ),
	.cout(Xd_0__inst_mult_13_473 ),
	.shareout(Xd_0__inst_mult_13_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_144 (
// Equation(s):
// Xd_0__inst_mult_13_476  = SUM(( (din_a[157] & din_b[165]) ) + ( Xd_0__inst_mult_13_462  ) + ( Xd_0__inst_mult_13_461  ))
// Xd_0__inst_mult_13_477  = CARRY(( (din_a[157] & din_b[165]) ) + ( Xd_0__inst_mult_13_462  ) + ( Xd_0__inst_mult_13_461  ))
// Xd_0__inst_mult_13_478  = SHARE((din_a[157] & din_b[166]))

	.dataa(!din_a[157]),
	.datab(!din_b[165]),
	.datac(!din_b[166]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_461 ),
	.sharein(Xd_0__inst_mult_13_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_476 ),
	.cout(Xd_0__inst_mult_13_477 ),
	.shareout(Xd_0__inst_mult_13_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_145 (
// Equation(s):
// Xd_0__inst_mult_13_480  = SUM(( (!din_a[159] & (((din_a[158] & din_b[164])))) # (din_a[159] & (!din_b[163] $ (((!din_a[158]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_586  ) + ( Xd_0__inst_mult_13_585  ))
// Xd_0__inst_mult_13_481  = CARRY(( (!din_a[159] & (((din_a[158] & din_b[164])))) # (din_a[159] & (!din_b[163] $ (((!din_a[158]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_586  ) + ( Xd_0__inst_mult_13_585  ))
// Xd_0__inst_mult_13_482  = SHARE((din_a[159] & (din_b[163] & (din_a[158] & din_b[164]))))

	.dataa(!din_a[159]),
	.datab(!din_b[163]),
	.datac(!din_a[158]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_585 ),
	.sharein(Xd_0__inst_mult_13_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_480 ),
	.cout(Xd_0__inst_mult_13_481 ),
	.shareout(Xd_0__inst_mult_13_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_145 (
// Equation(s):
// Xd_0__inst_mult_14_480  = SUM(( (din_a[173] & din_b[173]) ) + ( Xd_0__inst_mult_14_474  ) + ( Xd_0__inst_mult_14_473  ))
// Xd_0__inst_mult_14_481  = CARRY(( (din_a[173] & din_b[173]) ) + ( Xd_0__inst_mult_14_474  ) + ( Xd_0__inst_mult_14_473  ))
// Xd_0__inst_mult_14_482  = SHARE((din_a[173] & din_b[174]))

	.dataa(!din_a[173]),
	.datab(!din_b[173]),
	.datac(!din_b[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_473 ),
	.sharein(Xd_0__inst_mult_14_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_480 ),
	.cout(Xd_0__inst_mult_14_481 ),
	.shareout(Xd_0__inst_mult_14_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_146 (
// Equation(s):
// Xd_0__inst_mult_14_484  = SUM(( (din_a[169] & din_b[177]) ) + ( Xd_0__inst_mult_14_478  ) + ( Xd_0__inst_mult_14_477  ))
// Xd_0__inst_mult_14_485  = CARRY(( (din_a[169] & din_b[177]) ) + ( Xd_0__inst_mult_14_478  ) + ( Xd_0__inst_mult_14_477  ))
// Xd_0__inst_mult_14_486  = SHARE((din_a[169] & din_b[178]))

	.dataa(!din_a[169]),
	.datab(!din_b[177]),
	.datac(!din_b[178]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_477 ),
	.sharein(Xd_0__inst_mult_14_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_484 ),
	.cout(Xd_0__inst_mult_14_485 ),
	.shareout(Xd_0__inst_mult_14_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_147 (
// Equation(s):
// Xd_0__inst_mult_14_488  = SUM(( (!din_a[171] & (((din_a[170] & din_b[176])))) # (din_a[171] & (!din_b[175] $ (((!din_a[170]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_586  ) + ( Xd_0__inst_mult_14_585  ))
// Xd_0__inst_mult_14_489  = CARRY(( (!din_a[171] & (((din_a[170] & din_b[176])))) # (din_a[171] & (!din_b[175] $ (((!din_a[170]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_586  ) + ( Xd_0__inst_mult_14_585  ))
// Xd_0__inst_mult_14_490  = SHARE((din_a[171] & (din_b[175] & (din_a[170] & din_b[176]))))

	.dataa(!din_a[171]),
	.datab(!din_b[175]),
	.datac(!din_a[170]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_585 ),
	.sharein(Xd_0__inst_mult_14_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_488 ),
	.cout(Xd_0__inst_mult_14_489 ),
	.shareout(Xd_0__inst_mult_14_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_148 (
// Equation(s):
// Xd_0__inst_mult_15_492  = SUM(( (din_a[188] & din_b[182]) ) + ( Xd_0__inst_mult_15_478  ) + ( Xd_0__inst_mult_15_477  ))
// Xd_0__inst_mult_15_493  = CARRY(( (din_a[188] & din_b[182]) ) + ( Xd_0__inst_mult_15_478  ) + ( Xd_0__inst_mult_15_477  ))
// Xd_0__inst_mult_15_494  = SHARE((din_a[190] & din_b[181]))

	.dataa(!din_a[188]),
	.datab(!din_b[182]),
	.datac(!din_a[190]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_477 ),
	.sharein(Xd_0__inst_mult_15_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_492 ),
	.cout(Xd_0__inst_mult_15_493 ),
	.shareout(Xd_0__inst_mult_15_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_149 (
// Equation(s):
// Xd_0__inst_mult_15_496  = SUM(( (!din_a[187] & (((din_a[186] & din_b[184])))) # (din_a[187] & (!din_b[183] $ (((!din_a[186]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_482  ) + ( Xd_0__inst_mult_15_481  ))
// Xd_0__inst_mult_15_497  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[184])))) # (din_a[187] & (!din_b[183] $ (((!din_a[186]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_482  ) + ( Xd_0__inst_mult_15_481  ))
// Xd_0__inst_mult_15_498  = SHARE((din_a[187] & (din_b[183] & (din_a[186] & din_b[184]))))

	.dataa(!din_a[187]),
	.datab(!din_b[183]),
	.datac(!din_a[186]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_481 ),
	.sharein(Xd_0__inst_mult_15_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_496 ),
	.cout(Xd_0__inst_mult_15_497 ),
	.shareout(Xd_0__inst_mult_15_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_150 (
// Equation(s):
// Xd_0__inst_mult_15_500  = SUM(( (din_a[185] & din_b[185]) ) + ( Xd_0__inst_mult_15_486  ) + ( Xd_0__inst_mult_15_485  ))
// Xd_0__inst_mult_15_501  = CARRY(( (din_a[185] & din_b[185]) ) + ( Xd_0__inst_mult_15_486  ) + ( Xd_0__inst_mult_15_485  ))
// Xd_0__inst_mult_15_502  = SHARE((din_a[185] & din_b[186]))

	.dataa(!din_a[185]),
	.datab(!din_b[185]),
	.datac(!din_b[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_485 ),
	.sharein(Xd_0__inst_mult_15_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_500 ),
	.cout(Xd_0__inst_mult_15_501 ),
	.shareout(Xd_0__inst_mult_15_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_151 (
// Equation(s):
// Xd_0__inst_mult_15_504  = SUM(( (din_a[181] & din_b[189]) ) + ( Xd_0__inst_mult_15_490  ) + ( Xd_0__inst_mult_15_489  ))
// Xd_0__inst_mult_15_505  = CARRY(( (din_a[181] & din_b[189]) ) + ( Xd_0__inst_mult_15_490  ) + ( Xd_0__inst_mult_15_489  ))
// Xd_0__inst_mult_15_506  = SHARE((din_a[181] & din_b[190]))

	.dataa(!din_a[181]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_489 ),
	.sharein(Xd_0__inst_mult_15_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_504 ),
	.cout(Xd_0__inst_mult_15_505 ),
	.shareout(Xd_0__inst_mult_15_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_152 (
// Equation(s):
// Xd_0__inst_mult_15_508  = SUM(( (!din_a[183] & (((din_a[182] & din_b[188])))) # (din_a[183] & (!din_b[187] $ (((!din_a[182]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_582  ) + ( Xd_0__inst_mult_15_581  ))
// Xd_0__inst_mult_15_509  = CARRY(( (!din_a[183] & (((din_a[182] & din_b[188])))) # (din_a[183] & (!din_b[187] $ (((!din_a[182]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_582  ) + ( Xd_0__inst_mult_15_581  ))
// Xd_0__inst_mult_15_510  = SHARE((din_a[183] & (din_b[187] & (din_a[182] & din_b[188]))))

	.dataa(!din_a[183]),
	.datab(!din_b[187]),
	.datac(!din_a[182]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_581 ),
	.sharein(Xd_0__inst_mult_15_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_508 ),
	.cout(Xd_0__inst_mult_15_509 ),
	.shareout(Xd_0__inst_mult_15_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_137 (
// Equation(s):
// Xd_0__inst_mult_10_460  = SUM(( (din_a[128] & din_b[122]) ) + ( Xd_0__inst_mult_10_446  ) + ( Xd_0__inst_mult_10_445  ))
// Xd_0__inst_mult_10_461  = CARRY(( (din_a[128] & din_b[122]) ) + ( Xd_0__inst_mult_10_446  ) + ( Xd_0__inst_mult_10_445  ))
// Xd_0__inst_mult_10_462  = SHARE((din_a[130] & din_b[121]))

	.dataa(!din_a[128]),
	.datab(!din_b[122]),
	.datac(!din_a[130]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_445 ),
	.sharein(Xd_0__inst_mult_10_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_460 ),
	.cout(Xd_0__inst_mult_10_461 ),
	.shareout(Xd_0__inst_mult_10_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_138 (
// Equation(s):
// Xd_0__inst_mult_10_464  = SUM(( (!din_a[127] & (((din_a[126] & din_b[124])))) # (din_a[127] & (!din_b[123] $ (((!din_a[126]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_450  ) + ( Xd_0__inst_mult_10_449  ))
// Xd_0__inst_mult_10_465  = CARRY(( (!din_a[127] & (((din_a[126] & din_b[124])))) # (din_a[127] & (!din_b[123] $ (((!din_a[126]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_450  ) + ( Xd_0__inst_mult_10_449  ))
// Xd_0__inst_mult_10_466  = SHARE((din_a[127] & (din_b[123] & (din_a[126] & din_b[124]))))

	.dataa(!din_a[127]),
	.datab(!din_b[123]),
	.datac(!din_a[126]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_449 ),
	.sharein(Xd_0__inst_mult_10_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_464 ),
	.cout(Xd_0__inst_mult_10_465 ),
	.shareout(Xd_0__inst_mult_10_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_139 (
// Equation(s):
// Xd_0__inst_mult_10_468  = SUM(( (din_a[125] & din_b[125]) ) + ( Xd_0__inst_mult_10_454  ) + ( Xd_0__inst_mult_10_453  ))
// Xd_0__inst_mult_10_469  = CARRY(( (din_a[125] & din_b[125]) ) + ( Xd_0__inst_mult_10_454  ) + ( Xd_0__inst_mult_10_453  ))
// Xd_0__inst_mult_10_470  = SHARE((din_a[125] & din_b[126]))

	.dataa(!din_a[125]),
	.datab(!din_b[125]),
	.datac(!din_b[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_453 ),
	.sharein(Xd_0__inst_mult_10_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_468 ),
	.cout(Xd_0__inst_mult_10_469 ),
	.shareout(Xd_0__inst_mult_10_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_140 (
// Equation(s):
// Xd_0__inst_mult_10_472  = SUM(( (din_a[121] & din_b[129]) ) + ( Xd_0__inst_mult_10_458  ) + ( Xd_0__inst_mult_10_457  ))
// Xd_0__inst_mult_10_473  = CARRY(( (din_a[121] & din_b[129]) ) + ( Xd_0__inst_mult_10_458  ) + ( Xd_0__inst_mult_10_457  ))
// Xd_0__inst_mult_10_474  = SHARE((din_a[121] & din_b[130]))

	.dataa(!din_a[121]),
	.datab(!din_b[129]),
	.datac(!din_b[130]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_457 ),
	.sharein(Xd_0__inst_mult_10_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_472 ),
	.cout(Xd_0__inst_mult_10_473 ),
	.shareout(Xd_0__inst_mult_10_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_141 (
// Equation(s):
// Xd_0__inst_mult_10_476  = SUM(( (!din_a[123] & (((din_a[122] & din_b[128])))) # (din_a[123] & (!din_b[127] $ (((!din_a[122]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_582  ) + ( Xd_0__inst_mult_10_581  ))
// Xd_0__inst_mult_10_477  = CARRY(( (!din_a[123] & (((din_a[122] & din_b[128])))) # (din_a[123] & (!din_b[127] $ (((!din_a[122]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_582  ) + ( Xd_0__inst_mult_10_581  ))
// Xd_0__inst_mult_10_478  = SHARE((din_a[123] & (din_b[127] & (din_a[122] & din_b[128]))))

	.dataa(!din_a[123]),
	.datab(!din_b[127]),
	.datac(!din_a[122]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_581 ),
	.sharein(Xd_0__inst_mult_10_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_476 ),
	.cout(Xd_0__inst_mult_10_477 ),
	.shareout(Xd_0__inst_mult_10_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_141 (
// Equation(s):
// Xd_0__inst_mult_11_464  = SUM(( (din_a[140] & din_b[134]) ) + ( Xd_0__inst_mult_11_450  ) + ( Xd_0__inst_mult_11_449  ))
// Xd_0__inst_mult_11_465  = CARRY(( (din_a[140] & din_b[134]) ) + ( Xd_0__inst_mult_11_450  ) + ( Xd_0__inst_mult_11_449  ))
// Xd_0__inst_mult_11_466  = SHARE((din_a[142] & din_b[133]))

	.dataa(!din_a[140]),
	.datab(!din_b[134]),
	.datac(!din_a[142]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_449 ),
	.sharein(Xd_0__inst_mult_11_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_464 ),
	.cout(Xd_0__inst_mult_11_465 ),
	.shareout(Xd_0__inst_mult_11_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_142 (
// Equation(s):
// Xd_0__inst_mult_11_468  = SUM(( (!din_a[139] & (((din_a[138] & din_b[136])))) # (din_a[139] & (!din_b[135] $ (((!din_a[138]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_454  ) + ( Xd_0__inst_mult_11_453  ))
// Xd_0__inst_mult_11_469  = CARRY(( (!din_a[139] & (((din_a[138] & din_b[136])))) # (din_a[139] & (!din_b[135] $ (((!din_a[138]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_454  ) + ( Xd_0__inst_mult_11_453  ))
// Xd_0__inst_mult_11_470  = SHARE((din_a[139] & (din_b[135] & (din_a[138] & din_b[136]))))

	.dataa(!din_a[139]),
	.datab(!din_b[135]),
	.datac(!din_a[138]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_453 ),
	.sharein(Xd_0__inst_mult_11_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_468 ),
	.cout(Xd_0__inst_mult_11_469 ),
	.shareout(Xd_0__inst_mult_11_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_143 (
// Equation(s):
// Xd_0__inst_mult_11_472  = SUM(( (din_a[137] & din_b[137]) ) + ( Xd_0__inst_mult_11_458  ) + ( Xd_0__inst_mult_11_457  ))
// Xd_0__inst_mult_11_473  = CARRY(( (din_a[137] & din_b[137]) ) + ( Xd_0__inst_mult_11_458  ) + ( Xd_0__inst_mult_11_457  ))
// Xd_0__inst_mult_11_474  = SHARE((din_a[137] & din_b[138]))

	.dataa(!din_a[137]),
	.datab(!din_b[137]),
	.datac(!din_b[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_457 ),
	.sharein(Xd_0__inst_mult_11_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_472 ),
	.cout(Xd_0__inst_mult_11_473 ),
	.shareout(Xd_0__inst_mult_11_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_144 (
// Equation(s):
// Xd_0__inst_mult_11_476  = SUM(( (din_a[133] & din_b[141]) ) + ( Xd_0__inst_mult_11_462  ) + ( Xd_0__inst_mult_11_461  ))
// Xd_0__inst_mult_11_477  = CARRY(( (din_a[133] & din_b[141]) ) + ( Xd_0__inst_mult_11_462  ) + ( Xd_0__inst_mult_11_461  ))
// Xd_0__inst_mult_11_478  = SHARE((din_a[133] & din_b[142]))

	.dataa(!din_a[133]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_461 ),
	.sharein(Xd_0__inst_mult_11_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_476 ),
	.cout(Xd_0__inst_mult_11_477 ),
	.shareout(Xd_0__inst_mult_11_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_145 (
// Equation(s):
// Xd_0__inst_mult_11_480  = SUM(( (!din_a[135] & (((din_a[134] & din_b[140])))) # (din_a[135] & (!din_b[139] $ (((!din_a[134]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_586  ) + ( Xd_0__inst_mult_11_585  ))
// Xd_0__inst_mult_11_481  = CARRY(( (!din_a[135] & (((din_a[134] & din_b[140])))) # (din_a[135] & (!din_b[139] $ (((!din_a[134]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_586  ) + ( Xd_0__inst_mult_11_585  ))
// Xd_0__inst_mult_11_482  = SHARE((din_a[135] & (din_b[139] & (din_a[134] & din_b[140]))))

	.dataa(!din_a[135]),
	.datab(!din_b[139]),
	.datac(!din_a[134]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_585 ),
	.sharein(Xd_0__inst_mult_11_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_480 ),
	.cout(Xd_0__inst_mult_11_481 ),
	.shareout(Xd_0__inst_mult_11_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_141 (
// Equation(s):
// Xd_0__inst_mult_8_464  = SUM(( (din_a[104] & din_b[98]) ) + ( Xd_0__inst_mult_8_450  ) + ( Xd_0__inst_mult_8_449  ))
// Xd_0__inst_mult_8_465  = CARRY(( (din_a[104] & din_b[98]) ) + ( Xd_0__inst_mult_8_450  ) + ( Xd_0__inst_mult_8_449  ))
// Xd_0__inst_mult_8_466  = SHARE((din_a[106] & din_b[97]))

	.dataa(!din_a[104]),
	.datab(!din_b[98]),
	.datac(!din_a[106]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_449 ),
	.sharein(Xd_0__inst_mult_8_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_464 ),
	.cout(Xd_0__inst_mult_8_465 ),
	.shareout(Xd_0__inst_mult_8_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_142 (
// Equation(s):
// Xd_0__inst_mult_8_468  = SUM(( (!din_a[103] & (((din_a[102] & din_b[100])))) # (din_a[103] & (!din_b[99] $ (((!din_a[102]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_454  ) + ( Xd_0__inst_mult_8_453  ))
// Xd_0__inst_mult_8_469  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[100])))) # (din_a[103] & (!din_b[99] $ (((!din_a[102]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_454  ) + ( Xd_0__inst_mult_8_453  ))
// Xd_0__inst_mult_8_470  = SHARE((din_a[103] & (din_b[99] & (din_a[102] & din_b[100]))))

	.dataa(!din_a[103]),
	.datab(!din_b[99]),
	.datac(!din_a[102]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_453 ),
	.sharein(Xd_0__inst_mult_8_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_468 ),
	.cout(Xd_0__inst_mult_8_469 ),
	.shareout(Xd_0__inst_mult_8_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_143 (
// Equation(s):
// Xd_0__inst_mult_8_472  = SUM(( (din_a[101] & din_b[101]) ) + ( Xd_0__inst_mult_8_458  ) + ( Xd_0__inst_mult_8_457  ))
// Xd_0__inst_mult_8_473  = CARRY(( (din_a[101] & din_b[101]) ) + ( Xd_0__inst_mult_8_458  ) + ( Xd_0__inst_mult_8_457  ))
// Xd_0__inst_mult_8_474  = SHARE((din_a[101] & din_b[102]))

	.dataa(!din_a[101]),
	.datab(!din_b[101]),
	.datac(!din_b[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_457 ),
	.sharein(Xd_0__inst_mult_8_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_472 ),
	.cout(Xd_0__inst_mult_8_473 ),
	.shareout(Xd_0__inst_mult_8_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_144 (
// Equation(s):
// Xd_0__inst_mult_8_476  = SUM(( (din_a[97] & din_b[105]) ) + ( Xd_0__inst_mult_8_462  ) + ( Xd_0__inst_mult_8_461  ))
// Xd_0__inst_mult_8_477  = CARRY(( (din_a[97] & din_b[105]) ) + ( Xd_0__inst_mult_8_462  ) + ( Xd_0__inst_mult_8_461  ))
// Xd_0__inst_mult_8_478  = SHARE((din_a[97] & din_b[106]))

	.dataa(!din_a[97]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_461 ),
	.sharein(Xd_0__inst_mult_8_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_476 ),
	.cout(Xd_0__inst_mult_8_477 ),
	.shareout(Xd_0__inst_mult_8_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_145 (
// Equation(s):
// Xd_0__inst_mult_8_480  = SUM(( (!din_a[99] & (((din_a[98] & din_b[104])))) # (din_a[99] & (!din_b[103] $ (((!din_a[98]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_586  ) + ( Xd_0__inst_mult_8_585  ))
// Xd_0__inst_mult_8_481  = CARRY(( (!din_a[99] & (((din_a[98] & din_b[104])))) # (din_a[99] & (!din_b[103] $ (((!din_a[98]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_586  ) + ( Xd_0__inst_mult_8_585  ))
// Xd_0__inst_mult_8_482  = SHARE((din_a[99] & (din_b[103] & (din_a[98] & din_b[104]))))

	.dataa(!din_a[99]),
	.datab(!din_b[103]),
	.datac(!din_a[98]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_585 ),
	.sharein(Xd_0__inst_mult_8_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_480 ),
	.cout(Xd_0__inst_mult_8_481 ),
	.shareout(Xd_0__inst_mult_8_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_137 (
// Equation(s):
// Xd_0__inst_mult_9_460  = SUM(( (din_a[116] & din_b[110]) ) + ( Xd_0__inst_mult_9_446  ) + ( Xd_0__inst_mult_9_445  ))
// Xd_0__inst_mult_9_461  = CARRY(( (din_a[116] & din_b[110]) ) + ( Xd_0__inst_mult_9_446  ) + ( Xd_0__inst_mult_9_445  ))
// Xd_0__inst_mult_9_462  = SHARE((din_a[118] & din_b[109]))

	.dataa(!din_a[116]),
	.datab(!din_b[110]),
	.datac(!din_a[118]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_445 ),
	.sharein(Xd_0__inst_mult_9_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_460 ),
	.cout(Xd_0__inst_mult_9_461 ),
	.shareout(Xd_0__inst_mult_9_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_138 (
// Equation(s):
// Xd_0__inst_mult_9_464  = SUM(( (!din_a[115] & (((din_a[114] & din_b[112])))) # (din_a[115] & (!din_b[111] $ (((!din_a[114]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_450  ) + ( Xd_0__inst_mult_9_449  ))
// Xd_0__inst_mult_9_465  = CARRY(( (!din_a[115] & (((din_a[114] & din_b[112])))) # (din_a[115] & (!din_b[111] $ (((!din_a[114]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_450  ) + ( Xd_0__inst_mult_9_449  ))
// Xd_0__inst_mult_9_466  = SHARE((din_a[115] & (din_b[111] & (din_a[114] & din_b[112]))))

	.dataa(!din_a[115]),
	.datab(!din_b[111]),
	.datac(!din_a[114]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_449 ),
	.sharein(Xd_0__inst_mult_9_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_464 ),
	.cout(Xd_0__inst_mult_9_465 ),
	.shareout(Xd_0__inst_mult_9_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_139 (
// Equation(s):
// Xd_0__inst_mult_9_468  = SUM(( (din_a[113] & din_b[113]) ) + ( Xd_0__inst_mult_9_454  ) + ( Xd_0__inst_mult_9_453  ))
// Xd_0__inst_mult_9_469  = CARRY(( (din_a[113] & din_b[113]) ) + ( Xd_0__inst_mult_9_454  ) + ( Xd_0__inst_mult_9_453  ))
// Xd_0__inst_mult_9_470  = SHARE((din_a[113] & din_b[114]))

	.dataa(!din_a[113]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_453 ),
	.sharein(Xd_0__inst_mult_9_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_468 ),
	.cout(Xd_0__inst_mult_9_469 ),
	.shareout(Xd_0__inst_mult_9_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_140 (
// Equation(s):
// Xd_0__inst_mult_9_472  = SUM(( (din_a[109] & din_b[117]) ) + ( Xd_0__inst_mult_9_458  ) + ( Xd_0__inst_mult_9_457  ))
// Xd_0__inst_mult_9_473  = CARRY(( (din_a[109] & din_b[117]) ) + ( Xd_0__inst_mult_9_458  ) + ( Xd_0__inst_mult_9_457  ))
// Xd_0__inst_mult_9_474  = SHARE((din_a[109] & din_b[118]))

	.dataa(!din_a[109]),
	.datab(!din_b[117]),
	.datac(!din_b[118]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_457 ),
	.sharein(Xd_0__inst_mult_9_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_472 ),
	.cout(Xd_0__inst_mult_9_473 ),
	.shareout(Xd_0__inst_mult_9_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_141 (
// Equation(s):
// Xd_0__inst_mult_9_476  = SUM(( (!din_a[111] & (((din_a[110] & din_b[116])))) # (din_a[111] & (!din_b[115] $ (((!din_a[110]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_582  ) + ( Xd_0__inst_mult_9_581  ))
// Xd_0__inst_mult_9_477  = CARRY(( (!din_a[111] & (((din_a[110] & din_b[116])))) # (din_a[111] & (!din_b[115] $ (((!din_a[110]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_582  ) + ( Xd_0__inst_mult_9_581  ))
// Xd_0__inst_mult_9_478  = SHARE((din_a[111] & (din_b[115] & (din_a[110] & din_b[116]))))

	.dataa(!din_a[111]),
	.datab(!din_b[115]),
	.datac(!din_a[110]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_581 ),
	.sharein(Xd_0__inst_mult_9_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_476 ),
	.cout(Xd_0__inst_mult_9_477 ),
	.shareout(Xd_0__inst_mult_9_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_137 (
// Equation(s):
// Xd_0__inst_mult_6_460  = SUM(( (din_a[80] & din_b[74]) ) + ( Xd_0__inst_mult_6_446  ) + ( Xd_0__inst_mult_6_445  ))
// Xd_0__inst_mult_6_461  = CARRY(( (din_a[80] & din_b[74]) ) + ( Xd_0__inst_mult_6_446  ) + ( Xd_0__inst_mult_6_445  ))
// Xd_0__inst_mult_6_462  = SHARE((din_a[82] & din_b[73]))

	.dataa(!din_a[80]),
	.datab(!din_b[74]),
	.datac(!din_a[82]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_445 ),
	.sharein(Xd_0__inst_mult_6_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_460 ),
	.cout(Xd_0__inst_mult_6_461 ),
	.shareout(Xd_0__inst_mult_6_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_138 (
// Equation(s):
// Xd_0__inst_mult_6_464  = SUM(( (!din_a[79] & (((din_a[78] & din_b[76])))) # (din_a[79] & (!din_b[75] $ (((!din_a[78]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_450  ) + ( Xd_0__inst_mult_6_449  ))
// Xd_0__inst_mult_6_465  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[76])))) # (din_a[79] & (!din_b[75] $ (((!din_a[78]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_450  ) + ( Xd_0__inst_mult_6_449  ))
// Xd_0__inst_mult_6_466  = SHARE((din_a[79] & (din_b[75] & (din_a[78] & din_b[76]))))

	.dataa(!din_a[79]),
	.datab(!din_b[75]),
	.datac(!din_a[78]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_449 ),
	.sharein(Xd_0__inst_mult_6_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_464 ),
	.cout(Xd_0__inst_mult_6_465 ),
	.shareout(Xd_0__inst_mult_6_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_139 (
// Equation(s):
// Xd_0__inst_mult_6_468  = SUM(( (din_a[77] & din_b[77]) ) + ( Xd_0__inst_mult_6_454  ) + ( Xd_0__inst_mult_6_453  ))
// Xd_0__inst_mult_6_469  = CARRY(( (din_a[77] & din_b[77]) ) + ( Xd_0__inst_mult_6_454  ) + ( Xd_0__inst_mult_6_453  ))
// Xd_0__inst_mult_6_470  = SHARE((din_a[77] & din_b[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_453 ),
	.sharein(Xd_0__inst_mult_6_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_468 ),
	.cout(Xd_0__inst_mult_6_469 ),
	.shareout(Xd_0__inst_mult_6_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_140 (
// Equation(s):
// Xd_0__inst_mult_6_472  = SUM(( (din_a[73] & din_b[81]) ) + ( Xd_0__inst_mult_6_458  ) + ( Xd_0__inst_mult_6_457  ))
// Xd_0__inst_mult_6_473  = CARRY(( (din_a[73] & din_b[81]) ) + ( Xd_0__inst_mult_6_458  ) + ( Xd_0__inst_mult_6_457  ))
// Xd_0__inst_mult_6_474  = SHARE((din_a[73] & din_b[82]))

	.dataa(!din_a[73]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_457 ),
	.sharein(Xd_0__inst_mult_6_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_472 ),
	.cout(Xd_0__inst_mult_6_473 ),
	.shareout(Xd_0__inst_mult_6_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_141 (
// Equation(s):
// Xd_0__inst_mult_6_476  = SUM(( (!din_a[75] & (((din_a[74] & din_b[80])))) # (din_a[75] & (!din_b[79] $ (((!din_a[74]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_582  ) + ( Xd_0__inst_mult_6_581  ))
// Xd_0__inst_mult_6_477  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[80])))) # (din_a[75] & (!din_b[79] $ (((!din_a[74]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_582  ) + ( Xd_0__inst_mult_6_581  ))
// Xd_0__inst_mult_6_478  = SHARE((din_a[75] & (din_b[79] & (din_a[74] & din_b[80]))))

	.dataa(!din_a[75]),
	.datab(!din_b[79]),
	.datac(!din_a[74]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_581 ),
	.sharein(Xd_0__inst_mult_6_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_476 ),
	.cout(Xd_0__inst_mult_6_477 ),
	.shareout(Xd_0__inst_mult_6_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_133 (
// Equation(s):
// Xd_0__inst_mult_7_444  = SUM(( (din_a[92] & din_b[86]) ) + ( Xd_0__inst_mult_7_430  ) + ( Xd_0__inst_mult_7_429  ))
// Xd_0__inst_mult_7_445  = CARRY(( (din_a[92] & din_b[86]) ) + ( Xd_0__inst_mult_7_430  ) + ( Xd_0__inst_mult_7_429  ))
// Xd_0__inst_mult_7_446  = SHARE((din_a[94] & din_b[85]))

	.dataa(!din_a[92]),
	.datab(!din_b[86]),
	.datac(!din_a[94]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_429 ),
	.sharein(Xd_0__inst_mult_7_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_444 ),
	.cout(Xd_0__inst_mult_7_445 ),
	.shareout(Xd_0__inst_mult_7_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_134 (
// Equation(s):
// Xd_0__inst_mult_7_448  = SUM(( (!din_a[91] & (((din_a[90] & din_b[88])))) # (din_a[91] & (!din_b[87] $ (((!din_a[90]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_434  ) + ( Xd_0__inst_mult_7_433  ))
// Xd_0__inst_mult_7_449  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[88])))) # (din_a[91] & (!din_b[87] $ (((!din_a[90]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_434  ) + ( Xd_0__inst_mult_7_433  ))
// Xd_0__inst_mult_7_450  = SHARE((din_a[91] & (din_b[87] & (din_a[90] & din_b[88]))))

	.dataa(!din_a[91]),
	.datab(!din_b[87]),
	.datac(!din_a[90]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_433 ),
	.sharein(Xd_0__inst_mult_7_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_448 ),
	.cout(Xd_0__inst_mult_7_449 ),
	.shareout(Xd_0__inst_mult_7_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_135 (
// Equation(s):
// Xd_0__inst_mult_7_452  = SUM(( (din_a[89] & din_b[89]) ) + ( Xd_0__inst_mult_7_438  ) + ( Xd_0__inst_mult_7_437  ))
// Xd_0__inst_mult_7_453  = CARRY(( (din_a[89] & din_b[89]) ) + ( Xd_0__inst_mult_7_438  ) + ( Xd_0__inst_mult_7_437  ))
// Xd_0__inst_mult_7_454  = SHARE((din_a[89] & din_b[90]))

	.dataa(!din_a[89]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_437 ),
	.sharein(Xd_0__inst_mult_7_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_452 ),
	.cout(Xd_0__inst_mult_7_453 ),
	.shareout(Xd_0__inst_mult_7_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_136 (
// Equation(s):
// Xd_0__inst_mult_7_456  = SUM(( (din_a[85] & din_b[93]) ) + ( Xd_0__inst_mult_7_442  ) + ( Xd_0__inst_mult_7_441  ))
// Xd_0__inst_mult_7_457  = CARRY(( (din_a[85] & din_b[93]) ) + ( Xd_0__inst_mult_7_442  ) + ( Xd_0__inst_mult_7_441  ))
// Xd_0__inst_mult_7_458  = SHARE((din_a[85] & din_b[94]))

	.dataa(!din_a[85]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_441 ),
	.sharein(Xd_0__inst_mult_7_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_456 ),
	.cout(Xd_0__inst_mult_7_457 ),
	.shareout(Xd_0__inst_mult_7_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_137 (
// Equation(s):
// Xd_0__inst_mult_7_460  = SUM(( (!din_a[87] & (((din_a[86] & din_b[92])))) # (din_a[87] & (!din_b[91] $ (((!din_a[86]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_582  ) + ( Xd_0__inst_mult_7_581  ))
// Xd_0__inst_mult_7_461  = CARRY(( (!din_a[87] & (((din_a[86] & din_b[92])))) # (din_a[87] & (!din_b[91] $ (((!din_a[86]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_582  ) + ( Xd_0__inst_mult_7_581  ))
// Xd_0__inst_mult_7_462  = SHARE((din_a[87] & (din_b[91] & (din_a[86] & din_b[92]))))

	.dataa(!din_a[87]),
	.datab(!din_b[91]),
	.datac(!din_a[86]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_581 ),
	.sharein(Xd_0__inst_mult_7_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_460 ),
	.cout(Xd_0__inst_mult_7_461 ),
	.shareout(Xd_0__inst_mult_7_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_146 (
// Equation(s):
// Xd_0__inst_mult_4_484  = SUM(( (din_a[56] & din_b[50]) ) + ( Xd_0__inst_mult_4_470  ) + ( Xd_0__inst_mult_4_469  ))
// Xd_0__inst_mult_4_485  = CARRY(( (din_a[56] & din_b[50]) ) + ( Xd_0__inst_mult_4_470  ) + ( Xd_0__inst_mult_4_469  ))
// Xd_0__inst_mult_4_486  = SHARE((din_a[58] & din_b[49]))

	.dataa(!din_a[56]),
	.datab(!din_b[50]),
	.datac(!din_a[58]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_469 ),
	.sharein(Xd_0__inst_mult_4_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_484 ),
	.cout(Xd_0__inst_mult_4_485 ),
	.shareout(Xd_0__inst_mult_4_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_147 (
// Equation(s):
// Xd_0__inst_mult_4_488  = SUM(( (!din_a[55] & (((din_a[54] & din_b[52])))) # (din_a[55] & (!din_b[51] $ (((!din_a[54]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_474  ) + ( Xd_0__inst_mult_4_473  ))
// Xd_0__inst_mult_4_489  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[52])))) # (din_a[55] & (!din_b[51] $ (((!din_a[54]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_474  ) + ( Xd_0__inst_mult_4_473  ))
// Xd_0__inst_mult_4_490  = SHARE((din_a[55] & (din_b[51] & (din_a[54] & din_b[52]))))

	.dataa(!din_a[55]),
	.datab(!din_b[51]),
	.datac(!din_a[54]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_473 ),
	.sharein(Xd_0__inst_mult_4_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_488 ),
	.cout(Xd_0__inst_mult_4_489 ),
	.shareout(Xd_0__inst_mult_4_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_148 (
// Equation(s):
// Xd_0__inst_mult_4_492  = SUM(( (din_a[53] & din_b[53]) ) + ( Xd_0__inst_mult_4_478  ) + ( Xd_0__inst_mult_4_477  ))
// Xd_0__inst_mult_4_493  = CARRY(( (din_a[53] & din_b[53]) ) + ( Xd_0__inst_mult_4_478  ) + ( Xd_0__inst_mult_4_477  ))
// Xd_0__inst_mult_4_494  = SHARE((din_a[53] & din_b[54]))

	.dataa(!din_a[53]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_477 ),
	.sharein(Xd_0__inst_mult_4_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_492 ),
	.cout(Xd_0__inst_mult_4_493 ),
	.shareout(Xd_0__inst_mult_4_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_149 (
// Equation(s):
// Xd_0__inst_mult_4_496  = SUM(( (din_a[49] & din_b[57]) ) + ( Xd_0__inst_mult_4_482  ) + ( Xd_0__inst_mult_4_481  ))
// Xd_0__inst_mult_4_497  = CARRY(( (din_a[49] & din_b[57]) ) + ( Xd_0__inst_mult_4_482  ) + ( Xd_0__inst_mult_4_481  ))
// Xd_0__inst_mult_4_498  = SHARE((din_a[49] & din_b[58]))

	.dataa(!din_a[49]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_481 ),
	.sharein(Xd_0__inst_mult_4_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_496 ),
	.cout(Xd_0__inst_mult_4_497 ),
	.shareout(Xd_0__inst_mult_4_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_150 (
// Equation(s):
// Xd_0__inst_mult_4_500  = SUM(( (!din_a[51] & (((din_a[50] & din_b[56])))) # (din_a[51] & (!din_b[55] $ (((!din_a[50]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_582  ) + ( Xd_0__inst_mult_4_581  ))
// Xd_0__inst_mult_4_501  = CARRY(( (!din_a[51] & (((din_a[50] & din_b[56])))) # (din_a[51] & (!din_b[55] $ (((!din_a[50]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_582  ) + ( Xd_0__inst_mult_4_581  ))
// Xd_0__inst_mult_4_502  = SHARE((din_a[51] & (din_b[55] & (din_a[50] & din_b[56]))))

	.dataa(!din_a[51]),
	.datab(!din_b[55]),
	.datac(!din_a[50]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_581 ),
	.sharein(Xd_0__inst_mult_4_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_500 ),
	.cout(Xd_0__inst_mult_4_501 ),
	.shareout(Xd_0__inst_mult_4_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_133 (
// Equation(s):
// Xd_0__inst_mult_5_444  = SUM(( (din_a[68] & din_b[62]) ) + ( Xd_0__inst_mult_5_430  ) + ( Xd_0__inst_mult_5_429  ))
// Xd_0__inst_mult_5_445  = CARRY(( (din_a[68] & din_b[62]) ) + ( Xd_0__inst_mult_5_430  ) + ( Xd_0__inst_mult_5_429  ))
// Xd_0__inst_mult_5_446  = SHARE((din_a[70] & din_b[61]))

	.dataa(!din_a[68]),
	.datab(!din_b[62]),
	.datac(!din_a[70]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_429 ),
	.sharein(Xd_0__inst_mult_5_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_444 ),
	.cout(Xd_0__inst_mult_5_445 ),
	.shareout(Xd_0__inst_mult_5_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_134 (
// Equation(s):
// Xd_0__inst_mult_5_448  = SUM(( (!din_a[67] & (((din_a[66] & din_b[64])))) # (din_a[67] & (!din_b[63] $ (((!din_a[66]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_434  ) + ( Xd_0__inst_mult_5_433  ))
// Xd_0__inst_mult_5_449  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[64])))) # (din_a[67] & (!din_b[63] $ (((!din_a[66]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_434  ) + ( Xd_0__inst_mult_5_433  ))
// Xd_0__inst_mult_5_450  = SHARE((din_a[67] & (din_b[63] & (din_a[66] & din_b[64]))))

	.dataa(!din_a[67]),
	.datab(!din_b[63]),
	.datac(!din_a[66]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_433 ),
	.sharein(Xd_0__inst_mult_5_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_448 ),
	.cout(Xd_0__inst_mult_5_449 ),
	.shareout(Xd_0__inst_mult_5_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_135 (
// Equation(s):
// Xd_0__inst_mult_5_452  = SUM(( (din_a[65] & din_b[65]) ) + ( Xd_0__inst_mult_5_438  ) + ( Xd_0__inst_mult_5_437  ))
// Xd_0__inst_mult_5_453  = CARRY(( (din_a[65] & din_b[65]) ) + ( Xd_0__inst_mult_5_438  ) + ( Xd_0__inst_mult_5_437  ))
// Xd_0__inst_mult_5_454  = SHARE((din_a[65] & din_b[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_437 ),
	.sharein(Xd_0__inst_mult_5_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_452 ),
	.cout(Xd_0__inst_mult_5_453 ),
	.shareout(Xd_0__inst_mult_5_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_136 (
// Equation(s):
// Xd_0__inst_mult_5_456  = SUM(( (din_a[61] & din_b[69]) ) + ( Xd_0__inst_mult_5_442  ) + ( Xd_0__inst_mult_5_441  ))
// Xd_0__inst_mult_5_457  = CARRY(( (din_a[61] & din_b[69]) ) + ( Xd_0__inst_mult_5_442  ) + ( Xd_0__inst_mult_5_441  ))
// Xd_0__inst_mult_5_458  = SHARE((din_a[61] & din_b[70]))

	.dataa(!din_a[61]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_441 ),
	.sharein(Xd_0__inst_mult_5_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_456 ),
	.cout(Xd_0__inst_mult_5_457 ),
	.shareout(Xd_0__inst_mult_5_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_137 (
// Equation(s):
// Xd_0__inst_mult_5_460  = SUM(( (!din_a[63] & (((din_a[62] & din_b[68])))) # (din_a[63] & (!din_b[67] $ (((!din_a[62]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_582  ) + ( Xd_0__inst_mult_5_581  ))
// Xd_0__inst_mult_5_461  = CARRY(( (!din_a[63] & (((din_a[62] & din_b[68])))) # (din_a[63] & (!din_b[67] $ (((!din_a[62]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_582  ) + ( Xd_0__inst_mult_5_581  ))
// Xd_0__inst_mult_5_462  = SHARE((din_a[63] & (din_b[67] & (din_a[62] & din_b[68]))))

	.dataa(!din_a[63]),
	.datab(!din_b[67]),
	.datac(!din_a[62]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_581 ),
	.sharein(Xd_0__inst_mult_5_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_460 ),
	.cout(Xd_0__inst_mult_5_461 ),
	.shareout(Xd_0__inst_mult_5_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_137 (
// Equation(s):
// Xd_0__inst_mult_2_448  = SUM(( (din_a[32] & din_b[26]) ) + ( Xd_0__inst_mult_2_434  ) + ( Xd_0__inst_mult_2_433  ))
// Xd_0__inst_mult_2_449  = CARRY(( (din_a[32] & din_b[26]) ) + ( Xd_0__inst_mult_2_434  ) + ( Xd_0__inst_mult_2_433  ))
// Xd_0__inst_mult_2_450  = SHARE((din_a[34] & din_b[25]))

	.dataa(!din_a[32]),
	.datab(!din_b[26]),
	.datac(!din_a[34]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_433 ),
	.sharein(Xd_0__inst_mult_2_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_448 ),
	.cout(Xd_0__inst_mult_2_449 ),
	.shareout(Xd_0__inst_mult_2_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_138 (
// Equation(s):
// Xd_0__inst_mult_2_452  = SUM(( (!din_a[31] & (((din_a[30] & din_b[28])))) # (din_a[31] & (!din_b[27] $ (((!din_a[30]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_438  ) + ( Xd_0__inst_mult_2_437  ))
// Xd_0__inst_mult_2_453  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[28])))) # (din_a[31] & (!din_b[27] $ (((!din_a[30]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_438  ) + ( Xd_0__inst_mult_2_437  ))
// Xd_0__inst_mult_2_454  = SHARE((din_a[31] & (din_b[27] & (din_a[30] & din_b[28]))))

	.dataa(!din_a[31]),
	.datab(!din_b[27]),
	.datac(!din_a[30]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_437 ),
	.sharein(Xd_0__inst_mult_2_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_452 ),
	.cout(Xd_0__inst_mult_2_453 ),
	.shareout(Xd_0__inst_mult_2_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_67 (
// Equation(s):
// Xd_0__inst_mult_2_67_sumout  = SUM(( (din_a[34] & din_b[24]) ) + ( Xd_0__inst_mult_3_65  ) + ( Xd_0__inst_mult_3_64  ))
// Xd_0__inst_mult_2_68  = CARRY(( (din_a[34] & din_b[24]) ) + ( Xd_0__inst_mult_3_65  ) + ( Xd_0__inst_mult_3_64  ))
// Xd_0__inst_mult_2_69  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_64 ),
	.sharein(Xd_0__inst_mult_3_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_67_sumout ),
	.cout(Xd_0__inst_mult_2_68 ),
	.shareout(Xd_0__inst_mult_2_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_139 (
// Equation(s):
// Xd_0__inst_mult_2_456  = SUM(( (din_a[29] & din_b[29]) ) + ( Xd_0__inst_mult_2_442  ) + ( Xd_0__inst_mult_2_441  ))
// Xd_0__inst_mult_2_457  = CARRY(( (din_a[29] & din_b[29]) ) + ( Xd_0__inst_mult_2_442  ) + ( Xd_0__inst_mult_2_441  ))
// Xd_0__inst_mult_2_458  = SHARE((din_a[29] & din_b[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_441 ),
	.sharein(Xd_0__inst_mult_2_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_456 ),
	.cout(Xd_0__inst_mult_2_457 ),
	.shareout(Xd_0__inst_mult_2_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_140 (
// Equation(s):
// Xd_0__inst_mult_2_460  = SUM(( (din_a[25] & din_b[33]) ) + ( Xd_0__inst_mult_2_446  ) + ( Xd_0__inst_mult_2_445  ))
// Xd_0__inst_mult_2_461  = CARRY(( (din_a[25] & din_b[33]) ) + ( Xd_0__inst_mult_2_446  ) + ( Xd_0__inst_mult_2_445  ))
// Xd_0__inst_mult_2_462  = SHARE((din_a[25] & din_b[34]))

	.dataa(!din_a[25]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_445 ),
	.sharein(Xd_0__inst_mult_2_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_460 ),
	.cout(Xd_0__inst_mult_2_461 ),
	.shareout(Xd_0__inst_mult_2_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_141 (
// Equation(s):
// Xd_0__inst_mult_2_464  = SUM(( (!din_a[27] & (((din_a[26] & din_b[32])))) # (din_a[27] & (!din_b[31] $ (((!din_a[26]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_586  ) + ( Xd_0__inst_mult_2_585  ))
// Xd_0__inst_mult_2_465  = CARRY(( (!din_a[27] & (((din_a[26] & din_b[32])))) # (din_a[27] & (!din_b[31] $ (((!din_a[26]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_586  ) + ( Xd_0__inst_mult_2_585  ))
// Xd_0__inst_mult_2_466  = SHARE((din_a[27] & (din_b[31] & (din_a[26] & din_b[32]))))

	.dataa(!din_a[27]),
	.datab(!din_b[31]),
	.datac(!din_a[26]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_585 ),
	.sharein(Xd_0__inst_mult_2_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_464 ),
	.cout(Xd_0__inst_mult_2_465 ),
	.shareout(Xd_0__inst_mult_2_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_133 (
// Equation(s):
// Xd_0__inst_mult_3_444  = SUM(( (din_a[44] & din_b[38]) ) + ( Xd_0__inst_mult_3_430  ) + ( Xd_0__inst_mult_3_429  ))
// Xd_0__inst_mult_3_445  = CARRY(( (din_a[44] & din_b[38]) ) + ( Xd_0__inst_mult_3_430  ) + ( Xd_0__inst_mult_3_429  ))
// Xd_0__inst_mult_3_446  = SHARE((din_a[46] & din_b[37]))

	.dataa(!din_a[44]),
	.datab(!din_b[38]),
	.datac(!din_a[46]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_429 ),
	.sharein(Xd_0__inst_mult_3_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_444 ),
	.cout(Xd_0__inst_mult_3_445 ),
	.shareout(Xd_0__inst_mult_3_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_134 (
// Equation(s):
// Xd_0__inst_mult_3_448  = SUM(( (!din_a[43] & (((din_a[42] & din_b[40])))) # (din_a[43] & (!din_b[39] $ (((!din_a[42]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_434  ) + ( Xd_0__inst_mult_3_433  ))
// Xd_0__inst_mult_3_449  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[40])))) # (din_a[43] & (!din_b[39] $ (((!din_a[42]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_434  ) + ( Xd_0__inst_mult_3_433  ))
// Xd_0__inst_mult_3_450  = SHARE((din_a[43] & (din_b[39] & (din_a[42] & din_b[40]))))

	.dataa(!din_a[43]),
	.datab(!din_b[39]),
	.datac(!din_a[42]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_433 ),
	.sharein(Xd_0__inst_mult_3_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_448 ),
	.cout(Xd_0__inst_mult_3_449 ),
	.shareout(Xd_0__inst_mult_3_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_63 (
// Equation(s):
// Xd_0__inst_mult_3_63_sumout  = SUM(( (din_a[46] & din_b[36]) ) + ( Xd_0__inst_mult_0_69  ) + ( Xd_0__inst_mult_0_68  ))
// Xd_0__inst_mult_3_64  = CARRY(( (din_a[46] & din_b[36]) ) + ( Xd_0__inst_mult_0_69  ) + ( Xd_0__inst_mult_0_68  ))
// Xd_0__inst_mult_3_65  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_68 ),
	.sharein(Xd_0__inst_mult_0_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_63_sumout ),
	.cout(Xd_0__inst_mult_3_64 ),
	.shareout(Xd_0__inst_mult_3_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_135 (
// Equation(s):
// Xd_0__inst_mult_3_452  = SUM(( (din_a[41] & din_b[41]) ) + ( Xd_0__inst_mult_3_438  ) + ( Xd_0__inst_mult_3_437  ))
// Xd_0__inst_mult_3_453  = CARRY(( (din_a[41] & din_b[41]) ) + ( Xd_0__inst_mult_3_438  ) + ( Xd_0__inst_mult_3_437  ))
// Xd_0__inst_mult_3_454  = SHARE((din_a[41] & din_b[42]))

	.dataa(!din_a[41]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_437 ),
	.sharein(Xd_0__inst_mult_3_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_452 ),
	.cout(Xd_0__inst_mult_3_453 ),
	.shareout(Xd_0__inst_mult_3_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_136 (
// Equation(s):
// Xd_0__inst_mult_3_456  = SUM(( (din_a[37] & din_b[45]) ) + ( Xd_0__inst_mult_3_442  ) + ( Xd_0__inst_mult_3_441  ))
// Xd_0__inst_mult_3_457  = CARRY(( (din_a[37] & din_b[45]) ) + ( Xd_0__inst_mult_3_442  ) + ( Xd_0__inst_mult_3_441  ))
// Xd_0__inst_mult_3_458  = SHARE((din_a[37] & din_b[46]))

	.dataa(!din_a[37]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_441 ),
	.sharein(Xd_0__inst_mult_3_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_456 ),
	.cout(Xd_0__inst_mult_3_457 ),
	.shareout(Xd_0__inst_mult_3_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_137 (
// Equation(s):
// Xd_0__inst_mult_3_460  = SUM(( (!din_a[39] & (((din_a[38] & din_b[44])))) # (din_a[39] & (!din_b[43] $ (((!din_a[38]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_582  ) + ( Xd_0__inst_mult_3_581  ))
// Xd_0__inst_mult_3_461  = CARRY(( (!din_a[39] & (((din_a[38] & din_b[44])))) # (din_a[39] & (!din_b[43] $ (((!din_a[38]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_582  ) + ( Xd_0__inst_mult_3_581  ))
// Xd_0__inst_mult_3_462  = SHARE((din_a[39] & (din_b[43] & (din_a[38] & din_b[44]))))

	.dataa(!din_a[39]),
	.datab(!din_b[43]),
	.datac(!din_a[38]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_581 ),
	.sharein(Xd_0__inst_mult_3_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_460 ),
	.cout(Xd_0__inst_mult_3_461 ),
	.shareout(Xd_0__inst_mult_3_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_137 (
// Equation(s):
// Xd_0__inst_mult_0_448  = SUM(( (din_a[8] & din_b[2]) ) + ( Xd_0__inst_mult_0_434  ) + ( Xd_0__inst_mult_0_433  ))
// Xd_0__inst_mult_0_449  = CARRY(( (din_a[8] & din_b[2]) ) + ( Xd_0__inst_mult_0_434  ) + ( Xd_0__inst_mult_0_433  ))
// Xd_0__inst_mult_0_450  = SHARE((din_a[10] & din_b[1]))

	.dataa(!din_a[8]),
	.datab(!din_b[2]),
	.datac(!din_a[10]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_433 ),
	.sharein(Xd_0__inst_mult_0_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_448 ),
	.cout(Xd_0__inst_mult_0_449 ),
	.shareout(Xd_0__inst_mult_0_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_138 (
// Equation(s):
// Xd_0__inst_mult_0_452  = SUM(( (!din_a[7] & (((din_a[6] & din_b[4])))) # (din_a[7] & (!din_b[3] $ (((!din_a[6]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_438  ) + ( Xd_0__inst_mult_0_437  ))
// Xd_0__inst_mult_0_453  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[4])))) # (din_a[7] & (!din_b[3] $ (((!din_a[6]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_438  ) + ( Xd_0__inst_mult_0_437  ))
// Xd_0__inst_mult_0_454  = SHARE((din_a[7] & (din_b[3] & (din_a[6] & din_b[4]))))

	.dataa(!din_a[7]),
	.datab(!din_b[3]),
	.datac(!din_a[6]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_437 ),
	.sharein(Xd_0__inst_mult_0_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_452 ),
	.cout(Xd_0__inst_mult_0_453 ),
	.shareout(Xd_0__inst_mult_0_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_67 (
// Equation(s):
// Xd_0__inst_mult_0_67_sumout  = SUM(( (din_a[10] & din_b[0]) ) + ( Xd_0__inst_mult_15_69  ) + ( Xd_0__inst_mult_15_68  ))
// Xd_0__inst_mult_0_68  = CARRY(( (din_a[10] & din_b[0]) ) + ( Xd_0__inst_mult_15_69  ) + ( Xd_0__inst_mult_15_68  ))
// Xd_0__inst_mult_0_69  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_68 ),
	.sharein(Xd_0__inst_mult_15_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_67_sumout ),
	.cout(Xd_0__inst_mult_0_68 ),
	.shareout(Xd_0__inst_mult_0_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_139 (
// Equation(s):
// Xd_0__inst_mult_0_456  = SUM(( (din_a[5] & din_b[5]) ) + ( Xd_0__inst_mult_0_442  ) + ( Xd_0__inst_mult_0_441  ))
// Xd_0__inst_mult_0_457  = CARRY(( (din_a[5] & din_b[5]) ) + ( Xd_0__inst_mult_0_442  ) + ( Xd_0__inst_mult_0_441  ))
// Xd_0__inst_mult_0_458  = SHARE((din_a[5] & din_b[6]))

	.dataa(!din_a[5]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_441 ),
	.sharein(Xd_0__inst_mult_0_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_456 ),
	.cout(Xd_0__inst_mult_0_457 ),
	.shareout(Xd_0__inst_mult_0_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_140 (
// Equation(s):
// Xd_0__inst_mult_0_460  = SUM(( (din_a[1] & din_b[9]) ) + ( Xd_0__inst_mult_0_446  ) + ( Xd_0__inst_mult_0_445  ))
// Xd_0__inst_mult_0_461  = CARRY(( (din_a[1] & din_b[9]) ) + ( Xd_0__inst_mult_0_446  ) + ( Xd_0__inst_mult_0_445  ))
// Xd_0__inst_mult_0_462  = SHARE((din_a[1] & din_b[10]))

	.dataa(!din_a[1]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_445 ),
	.sharein(Xd_0__inst_mult_0_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_460 ),
	.cout(Xd_0__inst_mult_0_461 ),
	.shareout(Xd_0__inst_mult_0_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_141 (
// Equation(s):
// Xd_0__inst_mult_0_464  = SUM(( (!din_a[3] & (((din_a[2] & din_b[8])))) # (din_a[3] & (!din_b[7] $ (((!din_a[2]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_586  ) + ( Xd_0__inst_mult_0_585  ))
// Xd_0__inst_mult_0_465  = CARRY(( (!din_a[3] & (((din_a[2] & din_b[8])))) # (din_a[3] & (!din_b[7] $ (((!din_a[2]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_586  ) + ( Xd_0__inst_mult_0_585  ))
// Xd_0__inst_mult_0_466  = SHARE((din_a[3] & (din_b[7] & (din_a[2] & din_b[8]))))

	.dataa(!din_a[3]),
	.datab(!din_b[7]),
	.datac(!din_a[2]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_585 ),
	.sharein(Xd_0__inst_mult_0_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_464 ),
	.cout(Xd_0__inst_mult_0_465 ),
	.shareout(Xd_0__inst_mult_0_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_137 (
// Equation(s):
// Xd_0__inst_mult_1_448  = SUM(( (din_a[20] & din_b[14]) ) + ( Xd_0__inst_mult_1_434  ) + ( Xd_0__inst_mult_1_433  ))
// Xd_0__inst_mult_1_449  = CARRY(( (din_a[20] & din_b[14]) ) + ( Xd_0__inst_mult_1_434  ) + ( Xd_0__inst_mult_1_433  ))
// Xd_0__inst_mult_1_450  = SHARE((din_a[22] & din_b[13]))

	.dataa(!din_a[20]),
	.datab(!din_b[14]),
	.datac(!din_a[22]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_433 ),
	.sharein(Xd_0__inst_mult_1_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_448 ),
	.cout(Xd_0__inst_mult_1_449 ),
	.shareout(Xd_0__inst_mult_1_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_138 (
// Equation(s):
// Xd_0__inst_mult_1_452  = SUM(( (!din_a[19] & (((din_a[18] & din_b[16])))) # (din_a[19] & (!din_b[15] $ (((!din_a[18]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_438  ) + ( Xd_0__inst_mult_1_437  ))
// Xd_0__inst_mult_1_453  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[16])))) # (din_a[19] & (!din_b[15] $ (((!din_a[18]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_438  ) + ( Xd_0__inst_mult_1_437  ))
// Xd_0__inst_mult_1_454  = SHARE((din_a[19] & (din_b[15] & (din_a[18] & din_b[16]))))

	.dataa(!din_a[19]),
	.datab(!din_b[15]),
	.datac(!din_a[18]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_437 ),
	.sharein(Xd_0__inst_mult_1_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_452 ),
	.cout(Xd_0__inst_mult_1_453 ),
	.shareout(Xd_0__inst_mult_1_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_139 (
// Equation(s):
// Xd_0__inst_mult_1_456  = SUM(( (din_a[17] & din_b[17]) ) + ( Xd_0__inst_mult_1_442  ) + ( Xd_0__inst_mult_1_441  ))
// Xd_0__inst_mult_1_457  = CARRY(( (din_a[17] & din_b[17]) ) + ( Xd_0__inst_mult_1_442  ) + ( Xd_0__inst_mult_1_441  ))
// Xd_0__inst_mult_1_458  = SHARE((din_a[17] & din_b[18]))

	.dataa(!din_a[17]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_441 ),
	.sharein(Xd_0__inst_mult_1_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_456 ),
	.cout(Xd_0__inst_mult_1_457 ),
	.shareout(Xd_0__inst_mult_1_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_140 (
// Equation(s):
// Xd_0__inst_mult_1_460  = SUM(( (din_a[13] & din_b[21]) ) + ( Xd_0__inst_mult_1_446  ) + ( Xd_0__inst_mult_1_445  ))
// Xd_0__inst_mult_1_461  = CARRY(( (din_a[13] & din_b[21]) ) + ( Xd_0__inst_mult_1_446  ) + ( Xd_0__inst_mult_1_445  ))
// Xd_0__inst_mult_1_462  = SHARE((din_a[13] & din_b[22]))

	.dataa(!din_a[13]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_445 ),
	.sharein(Xd_0__inst_mult_1_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_460 ),
	.cout(Xd_0__inst_mult_1_461 ),
	.shareout(Xd_0__inst_mult_1_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_141 (
// Equation(s):
// Xd_0__inst_mult_1_464  = SUM(( (!din_a[15] & (((din_a[14] & din_b[20])))) # (din_a[15] & (!din_b[19] $ (((!din_a[14]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_586  ) + ( Xd_0__inst_mult_1_585  ))
// Xd_0__inst_mult_1_465  = CARRY(( (!din_a[15] & (((din_a[14] & din_b[20])))) # (din_a[15] & (!din_b[19] $ (((!din_a[14]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_586  ) + ( Xd_0__inst_mult_1_585  ))
// Xd_0__inst_mult_1_466  = SHARE((din_a[15] & (din_b[19] & (din_a[14] & din_b[20]))))

	.dataa(!din_a[15]),
	.datab(!din_b[19]),
	.datac(!din_a[14]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_585 ),
	.sharein(Xd_0__inst_mult_1_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_464 ),
	.cout(Xd_0__inst_mult_1_465 ),
	.shareout(Xd_0__inst_mult_1_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_149 (
// Equation(s):
// Xd_0__inst_mult_12_508  = SUM(( (din_a[153] & din_b[146]) ) + ( Xd_0__inst_mult_12_490  ) + ( Xd_0__inst_mult_12_489  ))
// Xd_0__inst_mult_12_509  = CARRY(( (din_a[153] & din_b[146]) ) + ( Xd_0__inst_mult_12_490  ) + ( Xd_0__inst_mult_12_489  ))
// Xd_0__inst_mult_12_510  = SHARE(GND)

	.dataa(!din_a[153]),
	.datab(!din_b[146]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_489 ),
	.sharein(Xd_0__inst_mult_12_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_508 ),
	.cout(Xd_0__inst_mult_12_509 ),
	.shareout(Xd_0__inst_mult_12_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_150 (
// Equation(s):
// Xd_0__inst_mult_12_512  = SUM(( (!din_a[152] & (((din_a[151] & din_b[148])))) # (din_a[152] & (!din_b[147] $ (((!din_a[151]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_494  ) + ( Xd_0__inst_mult_12_493  ))
// Xd_0__inst_mult_12_513  = CARRY(( (!din_a[152] & (((din_a[151] & din_b[148])))) # (din_a[152] & (!din_b[147] $ (((!din_a[151]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_12_494  ) + ( Xd_0__inst_mult_12_493  ))
// Xd_0__inst_mult_12_514  = SHARE((din_a[152] & (din_b[147] & (din_a[151] & din_b[148]))))

	.dataa(!din_a[152]),
	.datab(!din_b[147]),
	.datac(!din_a[151]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_493 ),
	.sharein(Xd_0__inst_mult_12_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_512 ),
	.cout(Xd_0__inst_mult_12_513 ),
	.shareout(Xd_0__inst_mult_12_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_151 (
// Equation(s):
// Xd_0__inst_mult_12_516  = SUM(( (din_a[150] & din_b[149]) ) + ( Xd_0__inst_mult_12_498  ) + ( Xd_0__inst_mult_12_497  ))
// Xd_0__inst_mult_12_517  = CARRY(( (din_a[150] & din_b[149]) ) + ( Xd_0__inst_mult_12_498  ) + ( Xd_0__inst_mult_12_497  ))
// Xd_0__inst_mult_12_518  = SHARE((din_a[150] & din_b[150]))

	.dataa(!din_a[150]),
	.datab(!din_b[149]),
	.datac(!din_b[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_497 ),
	.sharein(Xd_0__inst_mult_12_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_516 ),
	.cout(Xd_0__inst_mult_12_517 ),
	.shareout(Xd_0__inst_mult_12_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_152 (
// Equation(s):
// Xd_0__inst_mult_12_520  = SUM(( (din_a[146] & din_b[153]) ) + ( Xd_0__inst_mult_12_502  ) + ( Xd_0__inst_mult_12_501  ))
// Xd_0__inst_mult_12_521  = CARRY(( (din_a[146] & din_b[153]) ) + ( Xd_0__inst_mult_12_502  ) + ( Xd_0__inst_mult_12_501  ))
// Xd_0__inst_mult_12_522  = SHARE((din_a[146] & din_b[154]))

	.dataa(!din_a[146]),
	.datab(!din_b[153]),
	.datac(!din_b[154]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_501 ),
	.sharein(Xd_0__inst_mult_12_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_520 ),
	.cout(Xd_0__inst_mult_12_521 ),
	.shareout(Xd_0__inst_mult_12_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_153 (
// Equation(s):
// Xd_0__inst_mult_12_524  = SUM(( (!din_a[148] & (((din_a[147] & din_b[152])))) # (din_a[148] & (!din_b[151] $ (((!din_a[147]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_506  ) + ( Xd_0__inst_mult_12_505  ))
// Xd_0__inst_mult_12_525  = CARRY(( (!din_a[148] & (((din_a[147] & din_b[152])))) # (din_a[148] & (!din_b[151] $ (((!din_a[147]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_506  ) + ( Xd_0__inst_mult_12_505  ))
// Xd_0__inst_mult_12_526  = SHARE((din_a[148] & (din_b[151] & (din_a[147] & din_b[152]))))

	.dataa(!din_a[148]),
	.datab(!din_b[151]),
	.datac(!din_a[147]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_505 ),
	.sharein(Xd_0__inst_mult_12_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_524 ),
	.cout(Xd_0__inst_mult_12_525 ),
	.shareout(Xd_0__inst_mult_12_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_146 (
// Equation(s):
// Xd_0__inst_mult_13_484  = SUM(( (din_a[165] & din_b[158]) ) + ( Xd_0__inst_mult_13_466  ) + ( Xd_0__inst_mult_13_465  ))
// Xd_0__inst_mult_13_485  = CARRY(( (din_a[165] & din_b[158]) ) + ( Xd_0__inst_mult_13_466  ) + ( Xd_0__inst_mult_13_465  ))
// Xd_0__inst_mult_13_486  = SHARE(GND)

	.dataa(!din_a[165]),
	.datab(!din_b[158]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_465 ),
	.sharein(Xd_0__inst_mult_13_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_484 ),
	.cout(Xd_0__inst_mult_13_485 ),
	.shareout(Xd_0__inst_mult_13_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_147 (
// Equation(s):
// Xd_0__inst_mult_13_488  = SUM(( (!din_a[164] & (((din_a[163] & din_b[160])))) # (din_a[164] & (!din_b[159] $ (((!din_a[163]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_470  ) + ( Xd_0__inst_mult_13_469  ))
// Xd_0__inst_mult_13_489  = CARRY(( (!din_a[164] & (((din_a[163] & din_b[160])))) # (din_a[164] & (!din_b[159] $ (((!din_a[163]) # (!din_b[160]))))) ) + ( Xd_0__inst_mult_13_470  ) + ( Xd_0__inst_mult_13_469  ))
// Xd_0__inst_mult_13_490  = SHARE((din_a[164] & (din_b[159] & (din_a[163] & din_b[160]))))

	.dataa(!din_a[164]),
	.datab(!din_b[159]),
	.datac(!din_a[163]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_469 ),
	.sharein(Xd_0__inst_mult_13_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_488 ),
	.cout(Xd_0__inst_mult_13_489 ),
	.shareout(Xd_0__inst_mult_13_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_148 (
// Equation(s):
// Xd_0__inst_mult_13_492  = SUM(( (din_a[162] & din_b[161]) ) + ( Xd_0__inst_mult_13_474  ) + ( Xd_0__inst_mult_13_473  ))
// Xd_0__inst_mult_13_493  = CARRY(( (din_a[162] & din_b[161]) ) + ( Xd_0__inst_mult_13_474  ) + ( Xd_0__inst_mult_13_473  ))
// Xd_0__inst_mult_13_494  = SHARE((din_a[162] & din_b[162]))

	.dataa(!din_a[162]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_473 ),
	.sharein(Xd_0__inst_mult_13_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_492 ),
	.cout(Xd_0__inst_mult_13_493 ),
	.shareout(Xd_0__inst_mult_13_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_149 (
// Equation(s):
// Xd_0__inst_mult_13_496  = SUM(( (din_a[158] & din_b[165]) ) + ( Xd_0__inst_mult_13_478  ) + ( Xd_0__inst_mult_13_477  ))
// Xd_0__inst_mult_13_497  = CARRY(( (din_a[158] & din_b[165]) ) + ( Xd_0__inst_mult_13_478  ) + ( Xd_0__inst_mult_13_477  ))
// Xd_0__inst_mult_13_498  = SHARE((din_a[158] & din_b[166]))

	.dataa(!din_a[158]),
	.datab(!din_b[165]),
	.datac(!din_b[166]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_477 ),
	.sharein(Xd_0__inst_mult_13_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_496 ),
	.cout(Xd_0__inst_mult_13_497 ),
	.shareout(Xd_0__inst_mult_13_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_150 (
// Equation(s):
// Xd_0__inst_mult_13_500  = SUM(( (!din_a[160] & (((din_a[159] & din_b[164])))) # (din_a[160] & (!din_b[163] $ (((!din_a[159]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_482  ) + ( Xd_0__inst_mult_13_481  ))
// Xd_0__inst_mult_13_501  = CARRY(( (!din_a[160] & (((din_a[159] & din_b[164])))) # (din_a[160] & (!din_b[163] $ (((!din_a[159]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_482  ) + ( Xd_0__inst_mult_13_481  ))
// Xd_0__inst_mult_13_502  = SHARE((din_a[160] & (din_b[163] & (din_a[159] & din_b[164]))))

	.dataa(!din_a[160]),
	.datab(!din_b[163]),
	.datac(!din_a[159]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_481 ),
	.sharein(Xd_0__inst_mult_13_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_500 ),
	.cout(Xd_0__inst_mult_13_501 ),
	.shareout(Xd_0__inst_mult_13_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_148 (
// Equation(s):
// Xd_0__inst_mult_14_492  = SUM(( (din_a[174] & din_b[173]) ) + ( Xd_0__inst_mult_14_482  ) + ( Xd_0__inst_mult_14_481  ))
// Xd_0__inst_mult_14_493  = CARRY(( (din_a[174] & din_b[173]) ) + ( Xd_0__inst_mult_14_482  ) + ( Xd_0__inst_mult_14_481  ))
// Xd_0__inst_mult_14_494  = SHARE((din_a[174] & din_b[174]))

	.dataa(!din_a[174]),
	.datab(!din_b[173]),
	.datac(!din_b[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_481 ),
	.sharein(Xd_0__inst_mult_14_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_492 ),
	.cout(Xd_0__inst_mult_14_493 ),
	.shareout(Xd_0__inst_mult_14_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_149 (
// Equation(s):
// Xd_0__inst_mult_14_496  = SUM(( (din_a[170] & din_b[177]) ) + ( Xd_0__inst_mult_14_486  ) + ( Xd_0__inst_mult_14_485  ))
// Xd_0__inst_mult_14_497  = CARRY(( (din_a[170] & din_b[177]) ) + ( Xd_0__inst_mult_14_486  ) + ( Xd_0__inst_mult_14_485  ))
// Xd_0__inst_mult_14_498  = SHARE((din_a[170] & din_b[178]))

	.dataa(!din_a[170]),
	.datab(!din_b[177]),
	.datac(!din_b[178]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_485 ),
	.sharein(Xd_0__inst_mult_14_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_496 ),
	.cout(Xd_0__inst_mult_14_497 ),
	.shareout(Xd_0__inst_mult_14_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_150 (
// Equation(s):
// Xd_0__inst_mult_14_500  = SUM(( (!din_a[172] & (((din_a[171] & din_b[176])))) # (din_a[172] & (!din_b[175] $ (((!din_a[171]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_490  ) + ( Xd_0__inst_mult_14_489  ))
// Xd_0__inst_mult_14_501  = CARRY(( (!din_a[172] & (((din_a[171] & din_b[176])))) # (din_a[172] & (!din_b[175] $ (((!din_a[171]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_490  ) + ( Xd_0__inst_mult_14_489  ))
// Xd_0__inst_mult_14_502  = SHARE((din_a[172] & (din_b[175] & (din_a[171] & din_b[176]))))

	.dataa(!din_a[172]),
	.datab(!din_b[175]),
	.datac(!din_a[171]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_489 ),
	.sharein(Xd_0__inst_mult_14_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_500 ),
	.cout(Xd_0__inst_mult_14_501 ),
	.shareout(Xd_0__inst_mult_14_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_153 (
// Equation(s):
// Xd_0__inst_mult_15_512  = SUM(( (din_a[189] & din_b[182]) ) + ( Xd_0__inst_mult_15_494  ) + ( Xd_0__inst_mult_15_493  ))
// Xd_0__inst_mult_15_513  = CARRY(( (din_a[189] & din_b[182]) ) + ( Xd_0__inst_mult_15_494  ) + ( Xd_0__inst_mult_15_493  ))
// Xd_0__inst_mult_15_514  = SHARE(GND)

	.dataa(!din_a[189]),
	.datab(!din_b[182]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_493 ),
	.sharein(Xd_0__inst_mult_15_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_512 ),
	.cout(Xd_0__inst_mult_15_513 ),
	.shareout(Xd_0__inst_mult_15_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_154 (
// Equation(s):
// Xd_0__inst_mult_15_516  = SUM(( (!din_a[188] & (((din_a[187] & din_b[184])))) # (din_a[188] & (!din_b[183] $ (((!din_a[187]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_498  ) + ( Xd_0__inst_mult_15_497  ))
// Xd_0__inst_mult_15_517  = CARRY(( (!din_a[188] & (((din_a[187] & din_b[184])))) # (din_a[188] & (!din_b[183] $ (((!din_a[187]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_15_498  ) + ( Xd_0__inst_mult_15_497  ))
// Xd_0__inst_mult_15_518  = SHARE((din_a[188] & (din_b[183] & (din_a[187] & din_b[184]))))

	.dataa(!din_a[188]),
	.datab(!din_b[183]),
	.datac(!din_a[187]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_497 ),
	.sharein(Xd_0__inst_mult_15_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_516 ),
	.cout(Xd_0__inst_mult_15_517 ),
	.shareout(Xd_0__inst_mult_15_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_155 (
// Equation(s):
// Xd_0__inst_mult_15_520  = SUM(( (din_a[186] & din_b[185]) ) + ( Xd_0__inst_mult_15_502  ) + ( Xd_0__inst_mult_15_501  ))
// Xd_0__inst_mult_15_521  = CARRY(( (din_a[186] & din_b[185]) ) + ( Xd_0__inst_mult_15_502  ) + ( Xd_0__inst_mult_15_501  ))
// Xd_0__inst_mult_15_522  = SHARE((din_a[186] & din_b[186]))

	.dataa(!din_a[186]),
	.datab(!din_b[185]),
	.datac(!din_b[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_501 ),
	.sharein(Xd_0__inst_mult_15_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_520 ),
	.cout(Xd_0__inst_mult_15_521 ),
	.shareout(Xd_0__inst_mult_15_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_156 (
// Equation(s):
// Xd_0__inst_mult_15_524  = SUM(( (din_a[182] & din_b[189]) ) + ( Xd_0__inst_mult_15_506  ) + ( Xd_0__inst_mult_15_505  ))
// Xd_0__inst_mult_15_525  = CARRY(( (din_a[182] & din_b[189]) ) + ( Xd_0__inst_mult_15_506  ) + ( Xd_0__inst_mult_15_505  ))
// Xd_0__inst_mult_15_526  = SHARE((din_a[182] & din_b[190]))

	.dataa(!din_a[182]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_505 ),
	.sharein(Xd_0__inst_mult_15_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_524 ),
	.cout(Xd_0__inst_mult_15_525 ),
	.shareout(Xd_0__inst_mult_15_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_157 (
// Equation(s):
// Xd_0__inst_mult_15_528  = SUM(( (!din_a[184] & (((din_a[183] & din_b[188])))) # (din_a[184] & (!din_b[187] $ (((!din_a[183]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_510  ) + ( Xd_0__inst_mult_15_509  ))
// Xd_0__inst_mult_15_529  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[188])))) # (din_a[184] & (!din_b[187] $ (((!din_a[183]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_510  ) + ( Xd_0__inst_mult_15_509  ))
// Xd_0__inst_mult_15_530  = SHARE((din_a[184] & (din_b[187] & (din_a[183] & din_b[188]))))

	.dataa(!din_a[184]),
	.datab(!din_b[187]),
	.datac(!din_a[183]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_509 ),
	.sharein(Xd_0__inst_mult_15_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_528 ),
	.cout(Xd_0__inst_mult_15_529 ),
	.shareout(Xd_0__inst_mult_15_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_142 (
// Equation(s):
// Xd_0__inst_mult_10_480  = SUM(( (din_a[129] & din_b[122]) ) + ( Xd_0__inst_mult_10_462  ) + ( Xd_0__inst_mult_10_461  ))
// Xd_0__inst_mult_10_481  = CARRY(( (din_a[129] & din_b[122]) ) + ( Xd_0__inst_mult_10_462  ) + ( Xd_0__inst_mult_10_461  ))
// Xd_0__inst_mult_10_482  = SHARE(GND)

	.dataa(!din_a[129]),
	.datab(!din_b[122]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_461 ),
	.sharein(Xd_0__inst_mult_10_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_480 ),
	.cout(Xd_0__inst_mult_10_481 ),
	.shareout(Xd_0__inst_mult_10_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_143 (
// Equation(s):
// Xd_0__inst_mult_10_484  = SUM(( (!din_a[128] & (((din_a[127] & din_b[124])))) # (din_a[128] & (!din_b[123] $ (((!din_a[127]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_466  ) + ( Xd_0__inst_mult_10_465  ))
// Xd_0__inst_mult_10_485  = CARRY(( (!din_a[128] & (((din_a[127] & din_b[124])))) # (din_a[128] & (!din_b[123] $ (((!din_a[127]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_10_466  ) + ( Xd_0__inst_mult_10_465  ))
// Xd_0__inst_mult_10_486  = SHARE((din_a[128] & (din_b[123] & (din_a[127] & din_b[124]))))

	.dataa(!din_a[128]),
	.datab(!din_b[123]),
	.datac(!din_a[127]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_465 ),
	.sharein(Xd_0__inst_mult_10_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_484 ),
	.cout(Xd_0__inst_mult_10_485 ),
	.shareout(Xd_0__inst_mult_10_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_144 (
// Equation(s):
// Xd_0__inst_mult_10_488  = SUM(( (din_a[126] & din_b[125]) ) + ( Xd_0__inst_mult_10_470  ) + ( Xd_0__inst_mult_10_469  ))
// Xd_0__inst_mult_10_489  = CARRY(( (din_a[126] & din_b[125]) ) + ( Xd_0__inst_mult_10_470  ) + ( Xd_0__inst_mult_10_469  ))
// Xd_0__inst_mult_10_490  = SHARE((din_a[126] & din_b[126]))

	.dataa(!din_a[126]),
	.datab(!din_b[125]),
	.datac(!din_b[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_469 ),
	.sharein(Xd_0__inst_mult_10_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_488 ),
	.cout(Xd_0__inst_mult_10_489 ),
	.shareout(Xd_0__inst_mult_10_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_145 (
// Equation(s):
// Xd_0__inst_mult_10_492  = SUM(( (din_a[122] & din_b[129]) ) + ( Xd_0__inst_mult_10_474  ) + ( Xd_0__inst_mult_10_473  ))
// Xd_0__inst_mult_10_493  = CARRY(( (din_a[122] & din_b[129]) ) + ( Xd_0__inst_mult_10_474  ) + ( Xd_0__inst_mult_10_473  ))
// Xd_0__inst_mult_10_494  = SHARE((din_a[122] & din_b[130]))

	.dataa(!din_a[122]),
	.datab(!din_b[129]),
	.datac(!din_b[130]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_473 ),
	.sharein(Xd_0__inst_mult_10_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_492 ),
	.cout(Xd_0__inst_mult_10_493 ),
	.shareout(Xd_0__inst_mult_10_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_146 (
// Equation(s):
// Xd_0__inst_mult_10_496  = SUM(( (!din_a[124] & (((din_a[123] & din_b[128])))) # (din_a[124] & (!din_b[127] $ (((!din_a[123]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_478  ) + ( Xd_0__inst_mult_10_477  ))
// Xd_0__inst_mult_10_497  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[128])))) # (din_a[124] & (!din_b[127] $ (((!din_a[123]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_478  ) + ( Xd_0__inst_mult_10_477  ))
// Xd_0__inst_mult_10_498  = SHARE((din_a[124] & (din_b[127] & (din_a[123] & din_b[128]))))

	.dataa(!din_a[124]),
	.datab(!din_b[127]),
	.datac(!din_a[123]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_477 ),
	.sharein(Xd_0__inst_mult_10_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_496 ),
	.cout(Xd_0__inst_mult_10_497 ),
	.shareout(Xd_0__inst_mult_10_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_146 (
// Equation(s):
// Xd_0__inst_mult_11_484  = SUM(( (din_a[141] & din_b[134]) ) + ( Xd_0__inst_mult_11_466  ) + ( Xd_0__inst_mult_11_465  ))
// Xd_0__inst_mult_11_485  = CARRY(( (din_a[141] & din_b[134]) ) + ( Xd_0__inst_mult_11_466  ) + ( Xd_0__inst_mult_11_465  ))
// Xd_0__inst_mult_11_486  = SHARE(GND)

	.dataa(!din_a[141]),
	.datab(!din_b[134]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_465 ),
	.sharein(Xd_0__inst_mult_11_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_484 ),
	.cout(Xd_0__inst_mult_11_485 ),
	.shareout(Xd_0__inst_mult_11_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_147 (
// Equation(s):
// Xd_0__inst_mult_11_488  = SUM(( (!din_a[140] & (((din_a[139] & din_b[136])))) # (din_a[140] & (!din_b[135] $ (((!din_a[139]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_470  ) + ( Xd_0__inst_mult_11_469  ))
// Xd_0__inst_mult_11_489  = CARRY(( (!din_a[140] & (((din_a[139] & din_b[136])))) # (din_a[140] & (!din_b[135] $ (((!din_a[139]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_11_470  ) + ( Xd_0__inst_mult_11_469  ))
// Xd_0__inst_mult_11_490  = SHARE((din_a[140] & (din_b[135] & (din_a[139] & din_b[136]))))

	.dataa(!din_a[140]),
	.datab(!din_b[135]),
	.datac(!din_a[139]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_469 ),
	.sharein(Xd_0__inst_mult_11_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_488 ),
	.cout(Xd_0__inst_mult_11_489 ),
	.shareout(Xd_0__inst_mult_11_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_148 (
// Equation(s):
// Xd_0__inst_mult_11_492  = SUM(( (din_a[138] & din_b[137]) ) + ( Xd_0__inst_mult_11_474  ) + ( Xd_0__inst_mult_11_473  ))
// Xd_0__inst_mult_11_493  = CARRY(( (din_a[138] & din_b[137]) ) + ( Xd_0__inst_mult_11_474  ) + ( Xd_0__inst_mult_11_473  ))
// Xd_0__inst_mult_11_494  = SHARE((din_a[138] & din_b[138]))

	.dataa(!din_a[138]),
	.datab(!din_b[137]),
	.datac(!din_b[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_473 ),
	.sharein(Xd_0__inst_mult_11_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_492 ),
	.cout(Xd_0__inst_mult_11_493 ),
	.shareout(Xd_0__inst_mult_11_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_149 (
// Equation(s):
// Xd_0__inst_mult_11_496  = SUM(( (din_a[134] & din_b[141]) ) + ( Xd_0__inst_mult_11_478  ) + ( Xd_0__inst_mult_11_477  ))
// Xd_0__inst_mult_11_497  = CARRY(( (din_a[134] & din_b[141]) ) + ( Xd_0__inst_mult_11_478  ) + ( Xd_0__inst_mult_11_477  ))
// Xd_0__inst_mult_11_498  = SHARE((din_a[134] & din_b[142]))

	.dataa(!din_a[134]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_477 ),
	.sharein(Xd_0__inst_mult_11_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_496 ),
	.cout(Xd_0__inst_mult_11_497 ),
	.shareout(Xd_0__inst_mult_11_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_150 (
// Equation(s):
// Xd_0__inst_mult_11_500  = SUM(( (!din_a[136] & (((din_a[135] & din_b[140])))) # (din_a[136] & (!din_b[139] $ (((!din_a[135]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_482  ) + ( Xd_0__inst_mult_11_481  ))
// Xd_0__inst_mult_11_501  = CARRY(( (!din_a[136] & (((din_a[135] & din_b[140])))) # (din_a[136] & (!din_b[139] $ (((!din_a[135]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_482  ) + ( Xd_0__inst_mult_11_481  ))
// Xd_0__inst_mult_11_502  = SHARE((din_a[136] & (din_b[139] & (din_a[135] & din_b[140]))))

	.dataa(!din_a[136]),
	.datab(!din_b[139]),
	.datac(!din_a[135]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_481 ),
	.sharein(Xd_0__inst_mult_11_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_500 ),
	.cout(Xd_0__inst_mult_11_501 ),
	.shareout(Xd_0__inst_mult_11_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_146 (
// Equation(s):
// Xd_0__inst_mult_8_484  = SUM(( (din_a[105] & din_b[98]) ) + ( Xd_0__inst_mult_8_466  ) + ( Xd_0__inst_mult_8_465  ))
// Xd_0__inst_mult_8_485  = CARRY(( (din_a[105] & din_b[98]) ) + ( Xd_0__inst_mult_8_466  ) + ( Xd_0__inst_mult_8_465  ))
// Xd_0__inst_mult_8_486  = SHARE(GND)

	.dataa(!din_a[105]),
	.datab(!din_b[98]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_465 ),
	.sharein(Xd_0__inst_mult_8_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_484 ),
	.cout(Xd_0__inst_mult_8_485 ),
	.shareout(Xd_0__inst_mult_8_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_147 (
// Equation(s):
// Xd_0__inst_mult_8_488  = SUM(( (!din_a[104] & (((din_a[103] & din_b[100])))) # (din_a[104] & (!din_b[99] $ (((!din_a[103]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_470  ) + ( Xd_0__inst_mult_8_469  ))
// Xd_0__inst_mult_8_489  = CARRY(( (!din_a[104] & (((din_a[103] & din_b[100])))) # (din_a[104] & (!din_b[99] $ (((!din_a[103]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_8_470  ) + ( Xd_0__inst_mult_8_469  ))
// Xd_0__inst_mult_8_490  = SHARE((din_a[104] & (din_b[99] & (din_a[103] & din_b[100]))))

	.dataa(!din_a[104]),
	.datab(!din_b[99]),
	.datac(!din_a[103]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_469 ),
	.sharein(Xd_0__inst_mult_8_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_488 ),
	.cout(Xd_0__inst_mult_8_489 ),
	.shareout(Xd_0__inst_mult_8_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_148 (
// Equation(s):
// Xd_0__inst_mult_8_492  = SUM(( (din_a[102] & din_b[101]) ) + ( Xd_0__inst_mult_8_474  ) + ( Xd_0__inst_mult_8_473  ))
// Xd_0__inst_mult_8_493  = CARRY(( (din_a[102] & din_b[101]) ) + ( Xd_0__inst_mult_8_474  ) + ( Xd_0__inst_mult_8_473  ))
// Xd_0__inst_mult_8_494  = SHARE((din_a[102] & din_b[102]))

	.dataa(!din_a[102]),
	.datab(!din_b[101]),
	.datac(!din_b[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_473 ),
	.sharein(Xd_0__inst_mult_8_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_492 ),
	.cout(Xd_0__inst_mult_8_493 ),
	.shareout(Xd_0__inst_mult_8_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_149 (
// Equation(s):
// Xd_0__inst_mult_8_496  = SUM(( (din_a[98] & din_b[105]) ) + ( Xd_0__inst_mult_8_478  ) + ( Xd_0__inst_mult_8_477  ))
// Xd_0__inst_mult_8_497  = CARRY(( (din_a[98] & din_b[105]) ) + ( Xd_0__inst_mult_8_478  ) + ( Xd_0__inst_mult_8_477  ))
// Xd_0__inst_mult_8_498  = SHARE((din_a[98] & din_b[106]))

	.dataa(!din_a[98]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_477 ),
	.sharein(Xd_0__inst_mult_8_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_496 ),
	.cout(Xd_0__inst_mult_8_497 ),
	.shareout(Xd_0__inst_mult_8_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_150 (
// Equation(s):
// Xd_0__inst_mult_8_500  = SUM(( (!din_a[100] & (((din_a[99] & din_b[104])))) # (din_a[100] & (!din_b[103] $ (((!din_a[99]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_482  ) + ( Xd_0__inst_mult_8_481  ))
// Xd_0__inst_mult_8_501  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[104])))) # (din_a[100] & (!din_b[103] $ (((!din_a[99]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_482  ) + ( Xd_0__inst_mult_8_481  ))
// Xd_0__inst_mult_8_502  = SHARE((din_a[100] & (din_b[103] & (din_a[99] & din_b[104]))))

	.dataa(!din_a[100]),
	.datab(!din_b[103]),
	.datac(!din_a[99]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_481 ),
	.sharein(Xd_0__inst_mult_8_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_500 ),
	.cout(Xd_0__inst_mult_8_501 ),
	.shareout(Xd_0__inst_mult_8_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_142 (
// Equation(s):
// Xd_0__inst_mult_9_480  = SUM(( (din_a[117] & din_b[110]) ) + ( Xd_0__inst_mult_9_462  ) + ( Xd_0__inst_mult_9_461  ))
// Xd_0__inst_mult_9_481  = CARRY(( (din_a[117] & din_b[110]) ) + ( Xd_0__inst_mult_9_462  ) + ( Xd_0__inst_mult_9_461  ))
// Xd_0__inst_mult_9_482  = SHARE(GND)

	.dataa(!din_a[117]),
	.datab(!din_b[110]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_461 ),
	.sharein(Xd_0__inst_mult_9_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_480 ),
	.cout(Xd_0__inst_mult_9_481 ),
	.shareout(Xd_0__inst_mult_9_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_143 (
// Equation(s):
// Xd_0__inst_mult_9_484  = SUM(( (!din_a[116] & (((din_a[115] & din_b[112])))) # (din_a[116] & (!din_b[111] $ (((!din_a[115]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_466  ) + ( Xd_0__inst_mult_9_465  ))
// Xd_0__inst_mult_9_485  = CARRY(( (!din_a[116] & (((din_a[115] & din_b[112])))) # (din_a[116] & (!din_b[111] $ (((!din_a[115]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_9_466  ) + ( Xd_0__inst_mult_9_465  ))
// Xd_0__inst_mult_9_486  = SHARE((din_a[116] & (din_b[111] & (din_a[115] & din_b[112]))))

	.dataa(!din_a[116]),
	.datab(!din_b[111]),
	.datac(!din_a[115]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_465 ),
	.sharein(Xd_0__inst_mult_9_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_484 ),
	.cout(Xd_0__inst_mult_9_485 ),
	.shareout(Xd_0__inst_mult_9_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_144 (
// Equation(s):
// Xd_0__inst_mult_9_488  = SUM(( (din_a[114] & din_b[113]) ) + ( Xd_0__inst_mult_9_470  ) + ( Xd_0__inst_mult_9_469  ))
// Xd_0__inst_mult_9_489  = CARRY(( (din_a[114] & din_b[113]) ) + ( Xd_0__inst_mult_9_470  ) + ( Xd_0__inst_mult_9_469  ))
// Xd_0__inst_mult_9_490  = SHARE((din_a[114] & din_b[114]))

	.dataa(!din_a[114]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_469 ),
	.sharein(Xd_0__inst_mult_9_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_488 ),
	.cout(Xd_0__inst_mult_9_489 ),
	.shareout(Xd_0__inst_mult_9_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_145 (
// Equation(s):
// Xd_0__inst_mult_9_492  = SUM(( (din_a[110] & din_b[117]) ) + ( Xd_0__inst_mult_9_474  ) + ( Xd_0__inst_mult_9_473  ))
// Xd_0__inst_mult_9_493  = CARRY(( (din_a[110] & din_b[117]) ) + ( Xd_0__inst_mult_9_474  ) + ( Xd_0__inst_mult_9_473  ))
// Xd_0__inst_mult_9_494  = SHARE((din_a[110] & din_b[118]))

	.dataa(!din_a[110]),
	.datab(!din_b[117]),
	.datac(!din_b[118]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_473 ),
	.sharein(Xd_0__inst_mult_9_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_492 ),
	.cout(Xd_0__inst_mult_9_493 ),
	.shareout(Xd_0__inst_mult_9_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_146 (
// Equation(s):
// Xd_0__inst_mult_9_496  = SUM(( (!din_a[112] & (((din_a[111] & din_b[116])))) # (din_a[112] & (!din_b[115] $ (((!din_a[111]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_478  ) + ( Xd_0__inst_mult_9_477  ))
// Xd_0__inst_mult_9_497  = CARRY(( (!din_a[112] & (((din_a[111] & din_b[116])))) # (din_a[112] & (!din_b[115] $ (((!din_a[111]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_478  ) + ( Xd_0__inst_mult_9_477  ))
// Xd_0__inst_mult_9_498  = SHARE((din_a[112] & (din_b[115] & (din_a[111] & din_b[116]))))

	.dataa(!din_a[112]),
	.datab(!din_b[115]),
	.datac(!din_a[111]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_477 ),
	.sharein(Xd_0__inst_mult_9_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_496 ),
	.cout(Xd_0__inst_mult_9_497 ),
	.shareout(Xd_0__inst_mult_9_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_142 (
// Equation(s):
// Xd_0__inst_mult_6_480  = SUM(( (din_a[81] & din_b[74]) ) + ( Xd_0__inst_mult_6_462  ) + ( Xd_0__inst_mult_6_461  ))
// Xd_0__inst_mult_6_481  = CARRY(( (din_a[81] & din_b[74]) ) + ( Xd_0__inst_mult_6_462  ) + ( Xd_0__inst_mult_6_461  ))
// Xd_0__inst_mult_6_482  = SHARE(GND)

	.dataa(!din_a[81]),
	.datab(!din_b[74]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_461 ),
	.sharein(Xd_0__inst_mult_6_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_480 ),
	.cout(Xd_0__inst_mult_6_481 ),
	.shareout(Xd_0__inst_mult_6_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_143 (
// Equation(s):
// Xd_0__inst_mult_6_484  = SUM(( (!din_a[80] & (((din_a[79] & din_b[76])))) # (din_a[80] & (!din_b[75] $ (((!din_a[79]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_466  ) + ( Xd_0__inst_mult_6_465  ))
// Xd_0__inst_mult_6_485  = CARRY(( (!din_a[80] & (((din_a[79] & din_b[76])))) # (din_a[80] & (!din_b[75] $ (((!din_a[79]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_466  ) + ( Xd_0__inst_mult_6_465  ))
// Xd_0__inst_mult_6_486  = SHARE((din_a[80] & (din_b[75] & (din_a[79] & din_b[76]))))

	.dataa(!din_a[80]),
	.datab(!din_b[75]),
	.datac(!din_a[79]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_465 ),
	.sharein(Xd_0__inst_mult_6_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_484 ),
	.cout(Xd_0__inst_mult_6_485 ),
	.shareout(Xd_0__inst_mult_6_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_144 (
// Equation(s):
// Xd_0__inst_mult_6_488  = SUM(( (din_a[78] & din_b[77]) ) + ( Xd_0__inst_mult_6_470  ) + ( Xd_0__inst_mult_6_469  ))
// Xd_0__inst_mult_6_489  = CARRY(( (din_a[78] & din_b[77]) ) + ( Xd_0__inst_mult_6_470  ) + ( Xd_0__inst_mult_6_469  ))
// Xd_0__inst_mult_6_490  = SHARE((din_a[78] & din_b[78]))

	.dataa(!din_a[78]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_469 ),
	.sharein(Xd_0__inst_mult_6_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_488 ),
	.cout(Xd_0__inst_mult_6_489 ),
	.shareout(Xd_0__inst_mult_6_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_145 (
// Equation(s):
// Xd_0__inst_mult_6_492  = SUM(( (din_a[74] & din_b[81]) ) + ( Xd_0__inst_mult_6_474  ) + ( Xd_0__inst_mult_6_473  ))
// Xd_0__inst_mult_6_493  = CARRY(( (din_a[74] & din_b[81]) ) + ( Xd_0__inst_mult_6_474  ) + ( Xd_0__inst_mult_6_473  ))
// Xd_0__inst_mult_6_494  = SHARE((din_a[74] & din_b[82]))

	.dataa(!din_a[74]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_473 ),
	.sharein(Xd_0__inst_mult_6_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_492 ),
	.cout(Xd_0__inst_mult_6_493 ),
	.shareout(Xd_0__inst_mult_6_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_146 (
// Equation(s):
// Xd_0__inst_mult_6_496  = SUM(( (!din_a[76] & (((din_a[75] & din_b[80])))) # (din_a[76] & (!din_b[79] $ (((!din_a[75]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_478  ) + ( Xd_0__inst_mult_6_477  ))
// Xd_0__inst_mult_6_497  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[80])))) # (din_a[76] & (!din_b[79] $ (((!din_a[75]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_478  ) + ( Xd_0__inst_mult_6_477  ))
// Xd_0__inst_mult_6_498  = SHARE((din_a[76] & (din_b[79] & (din_a[75] & din_b[80]))))

	.dataa(!din_a[76]),
	.datab(!din_b[79]),
	.datac(!din_a[75]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_477 ),
	.sharein(Xd_0__inst_mult_6_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_496 ),
	.cout(Xd_0__inst_mult_6_497 ),
	.shareout(Xd_0__inst_mult_6_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_138 (
// Equation(s):
// Xd_0__inst_mult_7_464  = SUM(( (din_a[93] & din_b[86]) ) + ( Xd_0__inst_mult_7_446  ) + ( Xd_0__inst_mult_7_445  ))
// Xd_0__inst_mult_7_465  = CARRY(( (din_a[93] & din_b[86]) ) + ( Xd_0__inst_mult_7_446  ) + ( Xd_0__inst_mult_7_445  ))
// Xd_0__inst_mult_7_466  = SHARE(GND)

	.dataa(!din_a[93]),
	.datab(!din_b[86]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_445 ),
	.sharein(Xd_0__inst_mult_7_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_464 ),
	.cout(Xd_0__inst_mult_7_465 ),
	.shareout(Xd_0__inst_mult_7_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_139 (
// Equation(s):
// Xd_0__inst_mult_7_468  = SUM(( (!din_a[92] & (((din_a[91] & din_b[88])))) # (din_a[92] & (!din_b[87] $ (((!din_a[91]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_450  ) + ( Xd_0__inst_mult_7_449  ))
// Xd_0__inst_mult_7_469  = CARRY(( (!din_a[92] & (((din_a[91] & din_b[88])))) # (din_a[92] & (!din_b[87] $ (((!din_a[91]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_450  ) + ( Xd_0__inst_mult_7_449  ))
// Xd_0__inst_mult_7_470  = SHARE((din_a[92] & (din_b[87] & (din_a[91] & din_b[88]))))

	.dataa(!din_a[92]),
	.datab(!din_b[87]),
	.datac(!din_a[91]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_449 ),
	.sharein(Xd_0__inst_mult_7_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_468 ),
	.cout(Xd_0__inst_mult_7_469 ),
	.shareout(Xd_0__inst_mult_7_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_140 (
// Equation(s):
// Xd_0__inst_mult_7_472  = SUM(( (din_a[90] & din_b[89]) ) + ( Xd_0__inst_mult_7_454  ) + ( Xd_0__inst_mult_7_453  ))
// Xd_0__inst_mult_7_473  = CARRY(( (din_a[90] & din_b[89]) ) + ( Xd_0__inst_mult_7_454  ) + ( Xd_0__inst_mult_7_453  ))
// Xd_0__inst_mult_7_474  = SHARE((din_a[90] & din_b[90]))

	.dataa(!din_a[90]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_453 ),
	.sharein(Xd_0__inst_mult_7_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_472 ),
	.cout(Xd_0__inst_mult_7_473 ),
	.shareout(Xd_0__inst_mult_7_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_141 (
// Equation(s):
// Xd_0__inst_mult_7_476  = SUM(( (din_a[86] & din_b[93]) ) + ( Xd_0__inst_mult_7_458  ) + ( Xd_0__inst_mult_7_457  ))
// Xd_0__inst_mult_7_477  = CARRY(( (din_a[86] & din_b[93]) ) + ( Xd_0__inst_mult_7_458  ) + ( Xd_0__inst_mult_7_457  ))
// Xd_0__inst_mult_7_478  = SHARE((din_a[86] & din_b[94]))

	.dataa(!din_a[86]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_457 ),
	.sharein(Xd_0__inst_mult_7_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_476 ),
	.cout(Xd_0__inst_mult_7_477 ),
	.shareout(Xd_0__inst_mult_7_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_142 (
// Equation(s):
// Xd_0__inst_mult_7_480  = SUM(( (!din_a[88] & (((din_a[87] & din_b[92])))) # (din_a[88] & (!din_b[91] $ (((!din_a[87]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_462  ) + ( Xd_0__inst_mult_7_461  ))
// Xd_0__inst_mult_7_481  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[92])))) # (din_a[88] & (!din_b[91] $ (((!din_a[87]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_462  ) + ( Xd_0__inst_mult_7_461  ))
// Xd_0__inst_mult_7_482  = SHARE((din_a[88] & (din_b[91] & (din_a[87] & din_b[92]))))

	.dataa(!din_a[88]),
	.datab(!din_b[91]),
	.datac(!din_a[87]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_461 ),
	.sharein(Xd_0__inst_mult_7_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_480 ),
	.cout(Xd_0__inst_mult_7_481 ),
	.shareout(Xd_0__inst_mult_7_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_151 (
// Equation(s):
// Xd_0__inst_mult_4_504  = SUM(( (din_a[57] & din_b[50]) ) + ( Xd_0__inst_mult_4_486  ) + ( Xd_0__inst_mult_4_485  ))
// Xd_0__inst_mult_4_505  = CARRY(( (din_a[57] & din_b[50]) ) + ( Xd_0__inst_mult_4_486  ) + ( Xd_0__inst_mult_4_485  ))
// Xd_0__inst_mult_4_506  = SHARE(GND)

	.dataa(!din_a[57]),
	.datab(!din_b[50]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_485 ),
	.sharein(Xd_0__inst_mult_4_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_504 ),
	.cout(Xd_0__inst_mult_4_505 ),
	.shareout(Xd_0__inst_mult_4_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_152 (
// Equation(s):
// Xd_0__inst_mult_4_508  = SUM(( (!din_a[56] & (((din_a[55] & din_b[52])))) # (din_a[56] & (!din_b[51] $ (((!din_a[55]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_490  ) + ( Xd_0__inst_mult_4_489  ))
// Xd_0__inst_mult_4_509  = CARRY(( (!din_a[56] & (((din_a[55] & din_b[52])))) # (din_a[56] & (!din_b[51] $ (((!din_a[55]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_490  ) + ( Xd_0__inst_mult_4_489  ))
// Xd_0__inst_mult_4_510  = SHARE((din_a[56] & (din_b[51] & (din_a[55] & din_b[52]))))

	.dataa(!din_a[56]),
	.datab(!din_b[51]),
	.datac(!din_a[55]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_489 ),
	.sharein(Xd_0__inst_mult_4_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_508 ),
	.cout(Xd_0__inst_mult_4_509 ),
	.shareout(Xd_0__inst_mult_4_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_153 (
// Equation(s):
// Xd_0__inst_mult_4_512  = SUM(( (din_a[54] & din_b[53]) ) + ( Xd_0__inst_mult_4_494  ) + ( Xd_0__inst_mult_4_493  ))
// Xd_0__inst_mult_4_513  = CARRY(( (din_a[54] & din_b[53]) ) + ( Xd_0__inst_mult_4_494  ) + ( Xd_0__inst_mult_4_493  ))
// Xd_0__inst_mult_4_514  = SHARE((din_a[54] & din_b[54]))

	.dataa(!din_a[54]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_493 ),
	.sharein(Xd_0__inst_mult_4_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_512 ),
	.cout(Xd_0__inst_mult_4_513 ),
	.shareout(Xd_0__inst_mult_4_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_154 (
// Equation(s):
// Xd_0__inst_mult_4_516  = SUM(( (!din_a[52] & (((din_a[51] & din_b[56])))) # (din_a[52] & (!din_b[55] $ (((!din_a[51]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_502  ) + ( Xd_0__inst_mult_4_501  ))
// Xd_0__inst_mult_4_517  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[56])))) # (din_a[52] & (!din_b[55] $ (((!din_a[51]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_502  ) + ( Xd_0__inst_mult_4_501  ))
// Xd_0__inst_mult_4_518  = SHARE((din_a[52] & (din_b[55] & (din_a[51] & din_b[56]))))

	.dataa(!din_a[52]),
	.datab(!din_b[55]),
	.datac(!din_a[51]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_501 ),
	.sharein(Xd_0__inst_mult_4_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_516 ),
	.cout(Xd_0__inst_mult_4_517 ),
	.shareout(Xd_0__inst_mult_4_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_138 (
// Equation(s):
// Xd_0__inst_mult_5_464  = SUM(( (din_a[69] & din_b[62]) ) + ( Xd_0__inst_mult_5_446  ) + ( Xd_0__inst_mult_5_445  ))
// Xd_0__inst_mult_5_465  = CARRY(( (din_a[69] & din_b[62]) ) + ( Xd_0__inst_mult_5_446  ) + ( Xd_0__inst_mult_5_445  ))
// Xd_0__inst_mult_5_466  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[62]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_445 ),
	.sharein(Xd_0__inst_mult_5_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_464 ),
	.cout(Xd_0__inst_mult_5_465 ),
	.shareout(Xd_0__inst_mult_5_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_139 (
// Equation(s):
// Xd_0__inst_mult_5_468  = SUM(( (!din_a[68] & (((din_a[67] & din_b[64])))) # (din_a[68] & (!din_b[63] $ (((!din_a[67]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_450  ) + ( Xd_0__inst_mult_5_449  ))
// Xd_0__inst_mult_5_469  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[64])))) # (din_a[68] & (!din_b[63] $ (((!din_a[67]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_450  ) + ( Xd_0__inst_mult_5_449  ))
// Xd_0__inst_mult_5_470  = SHARE((din_a[68] & (din_b[63] & (din_a[67] & din_b[64]))))

	.dataa(!din_a[68]),
	.datab(!din_b[63]),
	.datac(!din_a[67]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_449 ),
	.sharein(Xd_0__inst_mult_5_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_468 ),
	.cout(Xd_0__inst_mult_5_469 ),
	.shareout(Xd_0__inst_mult_5_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_140 (
// Equation(s):
// Xd_0__inst_mult_5_472  = SUM(( (din_a[66] & din_b[65]) ) + ( Xd_0__inst_mult_5_454  ) + ( Xd_0__inst_mult_5_453  ))
// Xd_0__inst_mult_5_473  = CARRY(( (din_a[66] & din_b[65]) ) + ( Xd_0__inst_mult_5_454  ) + ( Xd_0__inst_mult_5_453  ))
// Xd_0__inst_mult_5_474  = SHARE((din_a[66] & din_b[66]))

	.dataa(!din_a[66]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_453 ),
	.sharein(Xd_0__inst_mult_5_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_472 ),
	.cout(Xd_0__inst_mult_5_473 ),
	.shareout(Xd_0__inst_mult_5_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_141 (
// Equation(s):
// Xd_0__inst_mult_5_476  = SUM(( (din_a[62] & din_b[69]) ) + ( Xd_0__inst_mult_5_458  ) + ( Xd_0__inst_mult_5_457  ))
// Xd_0__inst_mult_5_477  = CARRY(( (din_a[62] & din_b[69]) ) + ( Xd_0__inst_mult_5_458  ) + ( Xd_0__inst_mult_5_457  ))
// Xd_0__inst_mult_5_478  = SHARE((din_a[62] & din_b[70]))

	.dataa(!din_a[62]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_457 ),
	.sharein(Xd_0__inst_mult_5_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_476 ),
	.cout(Xd_0__inst_mult_5_477 ),
	.shareout(Xd_0__inst_mult_5_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_142 (
// Equation(s):
// Xd_0__inst_mult_5_480  = SUM(( (!din_a[64] & (((din_a[63] & din_b[68])))) # (din_a[64] & (!din_b[67] $ (((!din_a[63]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_462  ) + ( Xd_0__inst_mult_5_461  ))
// Xd_0__inst_mult_5_481  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[68])))) # (din_a[64] & (!din_b[67] $ (((!din_a[63]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_462  ) + ( Xd_0__inst_mult_5_461  ))
// Xd_0__inst_mult_5_482  = SHARE((din_a[64] & (din_b[67] & (din_a[63] & din_b[68]))))

	.dataa(!din_a[64]),
	.datab(!din_b[67]),
	.datac(!din_a[63]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_461 ),
	.sharein(Xd_0__inst_mult_5_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_480 ),
	.cout(Xd_0__inst_mult_5_481 ),
	.shareout(Xd_0__inst_mult_5_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_142 (
// Equation(s):
// Xd_0__inst_mult_2_468  = SUM(( (din_a[33] & din_b[26]) ) + ( Xd_0__inst_mult_2_450  ) + ( Xd_0__inst_mult_2_449  ))
// Xd_0__inst_mult_2_469  = CARRY(( (din_a[33] & din_b[26]) ) + ( Xd_0__inst_mult_2_450  ) + ( Xd_0__inst_mult_2_449  ))
// Xd_0__inst_mult_2_470  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[26]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_449 ),
	.sharein(Xd_0__inst_mult_2_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_468 ),
	.cout(Xd_0__inst_mult_2_469 ),
	.shareout(Xd_0__inst_mult_2_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_143 (
// Equation(s):
// Xd_0__inst_mult_2_472  = SUM(( (!din_a[32] & (((din_a[31] & din_b[28])))) # (din_a[32] & (!din_b[27] $ (((!din_a[31]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_454  ) + ( Xd_0__inst_mult_2_453  ))
// Xd_0__inst_mult_2_473  = CARRY(( (!din_a[32] & (((din_a[31] & din_b[28])))) # (din_a[32] & (!din_b[27] $ (((!din_a[31]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_454  ) + ( Xd_0__inst_mult_2_453  ))
// Xd_0__inst_mult_2_474  = SHARE((din_a[32] & (din_b[27] & (din_a[31] & din_b[28]))))

	.dataa(!din_a[32]),
	.datab(!din_b[27]),
	.datac(!din_a[31]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_453 ),
	.sharein(Xd_0__inst_mult_2_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_472 ),
	.cout(Xd_0__inst_mult_2_473 ),
	.shareout(Xd_0__inst_mult_2_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_144 (
// Equation(s):
// Xd_0__inst_mult_2_476  = SUM(( (din_a[30] & din_b[29]) ) + ( Xd_0__inst_mult_2_458  ) + ( Xd_0__inst_mult_2_457  ))
// Xd_0__inst_mult_2_477  = CARRY(( (din_a[30] & din_b[29]) ) + ( Xd_0__inst_mult_2_458  ) + ( Xd_0__inst_mult_2_457  ))
// Xd_0__inst_mult_2_478  = SHARE((din_a[30] & din_b[30]))

	.dataa(!din_a[30]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_457 ),
	.sharein(Xd_0__inst_mult_2_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_476 ),
	.cout(Xd_0__inst_mult_2_477 ),
	.shareout(Xd_0__inst_mult_2_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_145 (
// Equation(s):
// Xd_0__inst_mult_2_480  = SUM(( (din_a[26] & din_b[33]) ) + ( Xd_0__inst_mult_2_462  ) + ( Xd_0__inst_mult_2_461  ))
// Xd_0__inst_mult_2_481  = CARRY(( (din_a[26] & din_b[33]) ) + ( Xd_0__inst_mult_2_462  ) + ( Xd_0__inst_mult_2_461  ))
// Xd_0__inst_mult_2_482  = SHARE((din_a[26] & din_b[34]))

	.dataa(!din_a[26]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_461 ),
	.sharein(Xd_0__inst_mult_2_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_480 ),
	.cout(Xd_0__inst_mult_2_481 ),
	.shareout(Xd_0__inst_mult_2_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_146 (
// Equation(s):
// Xd_0__inst_mult_2_484  = SUM(( (!din_a[28] & (((din_a[27] & din_b[32])))) # (din_a[28] & (!din_b[31] $ (((!din_a[27]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_466  ) + ( Xd_0__inst_mult_2_465  ))
// Xd_0__inst_mult_2_485  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[32])))) # (din_a[28] & (!din_b[31] $ (((!din_a[27]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_466  ) + ( Xd_0__inst_mult_2_465  ))
// Xd_0__inst_mult_2_486  = SHARE((din_a[28] & (din_b[31] & (din_a[27] & din_b[32]))))

	.dataa(!din_a[28]),
	.datab(!din_b[31]),
	.datac(!din_a[27]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_465 ),
	.sharein(Xd_0__inst_mult_2_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_484 ),
	.cout(Xd_0__inst_mult_2_485 ),
	.shareout(Xd_0__inst_mult_2_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_138 (
// Equation(s):
// Xd_0__inst_mult_3_464  = SUM(( (din_a[45] & din_b[38]) ) + ( Xd_0__inst_mult_3_446  ) + ( Xd_0__inst_mult_3_445  ))
// Xd_0__inst_mult_3_465  = CARRY(( (din_a[45] & din_b[38]) ) + ( Xd_0__inst_mult_3_446  ) + ( Xd_0__inst_mult_3_445  ))
// Xd_0__inst_mult_3_466  = SHARE(GND)

	.dataa(!din_a[45]),
	.datab(!din_b[38]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_445 ),
	.sharein(Xd_0__inst_mult_3_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_464 ),
	.cout(Xd_0__inst_mult_3_465 ),
	.shareout(Xd_0__inst_mult_3_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_139 (
// Equation(s):
// Xd_0__inst_mult_3_468  = SUM(( (!din_a[44] & (((din_a[43] & din_b[40])))) # (din_a[44] & (!din_b[39] $ (((!din_a[43]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_450  ) + ( Xd_0__inst_mult_3_449  ))
// Xd_0__inst_mult_3_469  = CARRY(( (!din_a[44] & (((din_a[43] & din_b[40])))) # (din_a[44] & (!din_b[39] $ (((!din_a[43]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_450  ) + ( Xd_0__inst_mult_3_449  ))
// Xd_0__inst_mult_3_470  = SHARE((din_a[44] & (din_b[39] & (din_a[43] & din_b[40]))))

	.dataa(!din_a[44]),
	.datab(!din_b[39]),
	.datac(!din_a[43]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_449 ),
	.sharein(Xd_0__inst_mult_3_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_468 ),
	.cout(Xd_0__inst_mult_3_469 ),
	.shareout(Xd_0__inst_mult_3_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_140 (
// Equation(s):
// Xd_0__inst_mult_3_472  = SUM(( (din_a[42] & din_b[41]) ) + ( Xd_0__inst_mult_3_454  ) + ( Xd_0__inst_mult_3_453  ))
// Xd_0__inst_mult_3_473  = CARRY(( (din_a[42] & din_b[41]) ) + ( Xd_0__inst_mult_3_454  ) + ( Xd_0__inst_mult_3_453  ))
// Xd_0__inst_mult_3_474  = SHARE((din_a[42] & din_b[42]))

	.dataa(!din_a[42]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_453 ),
	.sharein(Xd_0__inst_mult_3_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_472 ),
	.cout(Xd_0__inst_mult_3_473 ),
	.shareout(Xd_0__inst_mult_3_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_141 (
// Equation(s):
// Xd_0__inst_mult_3_476  = SUM(( (din_a[38] & din_b[45]) ) + ( Xd_0__inst_mult_3_458  ) + ( Xd_0__inst_mult_3_457  ))
// Xd_0__inst_mult_3_477  = CARRY(( (din_a[38] & din_b[45]) ) + ( Xd_0__inst_mult_3_458  ) + ( Xd_0__inst_mult_3_457  ))
// Xd_0__inst_mult_3_478  = SHARE((din_a[38] & din_b[46]))

	.dataa(!din_a[38]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_457 ),
	.sharein(Xd_0__inst_mult_3_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_476 ),
	.cout(Xd_0__inst_mult_3_477 ),
	.shareout(Xd_0__inst_mult_3_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_142 (
// Equation(s):
// Xd_0__inst_mult_3_480  = SUM(( (!din_a[40] & (((din_a[39] & din_b[44])))) # (din_a[40] & (!din_b[43] $ (((!din_a[39]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_462  ) + ( Xd_0__inst_mult_3_461  ))
// Xd_0__inst_mult_3_481  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[44])))) # (din_a[40] & (!din_b[43] $ (((!din_a[39]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_462  ) + ( Xd_0__inst_mult_3_461  ))
// Xd_0__inst_mult_3_482  = SHARE((din_a[40] & (din_b[43] & (din_a[39] & din_b[44]))))

	.dataa(!din_a[40]),
	.datab(!din_b[43]),
	.datac(!din_a[39]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_461 ),
	.sharein(Xd_0__inst_mult_3_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_480 ),
	.cout(Xd_0__inst_mult_3_481 ),
	.shareout(Xd_0__inst_mult_3_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_142 (
// Equation(s):
// Xd_0__inst_mult_0_468  = SUM(( (din_a[9] & din_b[2]) ) + ( Xd_0__inst_mult_0_450  ) + ( Xd_0__inst_mult_0_449  ))
// Xd_0__inst_mult_0_469  = CARRY(( (din_a[9] & din_b[2]) ) + ( Xd_0__inst_mult_0_450  ) + ( Xd_0__inst_mult_0_449  ))
// Xd_0__inst_mult_0_470  = SHARE(GND)

	.dataa(!din_a[9]),
	.datab(!din_b[2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_449 ),
	.sharein(Xd_0__inst_mult_0_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_468 ),
	.cout(Xd_0__inst_mult_0_469 ),
	.shareout(Xd_0__inst_mult_0_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_143 (
// Equation(s):
// Xd_0__inst_mult_0_472  = SUM(( (!din_a[8] & (((din_a[7] & din_b[4])))) # (din_a[8] & (!din_b[3] $ (((!din_a[7]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_454  ) + ( Xd_0__inst_mult_0_453  ))
// Xd_0__inst_mult_0_473  = CARRY(( (!din_a[8] & (((din_a[7] & din_b[4])))) # (din_a[8] & (!din_b[3] $ (((!din_a[7]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_454  ) + ( Xd_0__inst_mult_0_453  ))
// Xd_0__inst_mult_0_474  = SHARE((din_a[8] & (din_b[3] & (din_a[7] & din_b[4]))))

	.dataa(!din_a[8]),
	.datab(!din_b[3]),
	.datac(!din_a[7]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_453 ),
	.sharein(Xd_0__inst_mult_0_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_472 ),
	.cout(Xd_0__inst_mult_0_473 ),
	.shareout(Xd_0__inst_mult_0_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_144 (
// Equation(s):
// Xd_0__inst_mult_0_476  = SUM(( (din_a[6] & din_b[5]) ) + ( Xd_0__inst_mult_0_458  ) + ( Xd_0__inst_mult_0_457  ))
// Xd_0__inst_mult_0_477  = CARRY(( (din_a[6] & din_b[5]) ) + ( Xd_0__inst_mult_0_458  ) + ( Xd_0__inst_mult_0_457  ))
// Xd_0__inst_mult_0_478  = SHARE((din_a[6] & din_b[6]))

	.dataa(!din_a[6]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_457 ),
	.sharein(Xd_0__inst_mult_0_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_476 ),
	.cout(Xd_0__inst_mult_0_477 ),
	.shareout(Xd_0__inst_mult_0_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_145 (
// Equation(s):
// Xd_0__inst_mult_0_480  = SUM(( (din_a[2] & din_b[9]) ) + ( Xd_0__inst_mult_0_462  ) + ( Xd_0__inst_mult_0_461  ))
// Xd_0__inst_mult_0_481  = CARRY(( (din_a[2] & din_b[9]) ) + ( Xd_0__inst_mult_0_462  ) + ( Xd_0__inst_mult_0_461  ))
// Xd_0__inst_mult_0_482  = SHARE((din_a[2] & din_b[10]))

	.dataa(!din_a[2]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_461 ),
	.sharein(Xd_0__inst_mult_0_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_480 ),
	.cout(Xd_0__inst_mult_0_481 ),
	.shareout(Xd_0__inst_mult_0_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_146 (
// Equation(s):
// Xd_0__inst_mult_0_484  = SUM(( (!din_a[4] & (((din_a[3] & din_b[8])))) # (din_a[4] & (!din_b[7] $ (((!din_a[3]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_466  ) + ( Xd_0__inst_mult_0_465  ))
// Xd_0__inst_mult_0_485  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[8])))) # (din_a[4] & (!din_b[7] $ (((!din_a[3]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_466  ) + ( Xd_0__inst_mult_0_465  ))
// Xd_0__inst_mult_0_486  = SHARE((din_a[4] & (din_b[7] & (din_a[3] & din_b[8]))))

	.dataa(!din_a[4]),
	.datab(!din_b[7]),
	.datac(!din_a[3]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_465 ),
	.sharein(Xd_0__inst_mult_0_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_484 ),
	.cout(Xd_0__inst_mult_0_485 ),
	.shareout(Xd_0__inst_mult_0_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_142 (
// Equation(s):
// Xd_0__inst_mult_1_468  = SUM(( (din_a[21] & din_b[14]) ) + ( Xd_0__inst_mult_1_450  ) + ( Xd_0__inst_mult_1_449  ))
// Xd_0__inst_mult_1_469  = CARRY(( (din_a[21] & din_b[14]) ) + ( Xd_0__inst_mult_1_450  ) + ( Xd_0__inst_mult_1_449  ))
// Xd_0__inst_mult_1_470  = SHARE(GND)

	.dataa(!din_a[21]),
	.datab(!din_b[14]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_449 ),
	.sharein(Xd_0__inst_mult_1_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_468 ),
	.cout(Xd_0__inst_mult_1_469 ),
	.shareout(Xd_0__inst_mult_1_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_143 (
// Equation(s):
// Xd_0__inst_mult_1_472  = SUM(( (!din_a[20] & (((din_a[19] & din_b[16])))) # (din_a[20] & (!din_b[15] $ (((!din_a[19]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_454  ) + ( Xd_0__inst_mult_1_453  ))
// Xd_0__inst_mult_1_473  = CARRY(( (!din_a[20] & (((din_a[19] & din_b[16])))) # (din_a[20] & (!din_b[15] $ (((!din_a[19]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_454  ) + ( Xd_0__inst_mult_1_453  ))
// Xd_0__inst_mult_1_474  = SHARE((din_a[20] & (din_b[15] & (din_a[19] & din_b[16]))))

	.dataa(!din_a[20]),
	.datab(!din_b[15]),
	.datac(!din_a[19]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_453 ),
	.sharein(Xd_0__inst_mult_1_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_472 ),
	.cout(Xd_0__inst_mult_1_473 ),
	.shareout(Xd_0__inst_mult_1_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_144 (
// Equation(s):
// Xd_0__inst_mult_1_476  = SUM(( (din_a[18] & din_b[17]) ) + ( Xd_0__inst_mult_1_458  ) + ( Xd_0__inst_mult_1_457  ))
// Xd_0__inst_mult_1_477  = CARRY(( (din_a[18] & din_b[17]) ) + ( Xd_0__inst_mult_1_458  ) + ( Xd_0__inst_mult_1_457  ))
// Xd_0__inst_mult_1_478  = SHARE((din_a[18] & din_b[18]))

	.dataa(!din_a[18]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_457 ),
	.sharein(Xd_0__inst_mult_1_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_476 ),
	.cout(Xd_0__inst_mult_1_477 ),
	.shareout(Xd_0__inst_mult_1_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_145 (
// Equation(s):
// Xd_0__inst_mult_1_480  = SUM(( (din_a[14] & din_b[21]) ) + ( Xd_0__inst_mult_1_462  ) + ( Xd_0__inst_mult_1_461  ))
// Xd_0__inst_mult_1_481  = CARRY(( (din_a[14] & din_b[21]) ) + ( Xd_0__inst_mult_1_462  ) + ( Xd_0__inst_mult_1_461  ))
// Xd_0__inst_mult_1_482  = SHARE((din_a[14] & din_b[22]))

	.dataa(!din_a[14]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_461 ),
	.sharein(Xd_0__inst_mult_1_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_480 ),
	.cout(Xd_0__inst_mult_1_481 ),
	.shareout(Xd_0__inst_mult_1_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_146 (
// Equation(s):
// Xd_0__inst_mult_1_484  = SUM(( (!din_a[16] & (((din_a[15] & din_b[20])))) # (din_a[16] & (!din_b[19] $ (((!din_a[15]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_466  ) + ( Xd_0__inst_mult_1_465  ))
// Xd_0__inst_mult_1_485  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[20])))) # (din_a[16] & (!din_b[19] $ (((!din_a[15]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_466  ) + ( Xd_0__inst_mult_1_465  ))
// Xd_0__inst_mult_1_486  = SHARE((din_a[16] & (din_b[19] & (din_a[15] & din_b[20]))))

	.dataa(!din_a[16]),
	.datab(!din_b[19]),
	.datac(!din_a[15]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_465 ),
	.sharein(Xd_0__inst_mult_1_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_484 ),
	.cout(Xd_0__inst_mult_1_485 ),
	.shareout(Xd_0__inst_mult_1_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_154 (
// Equation(s):
// Xd_0__inst_mult_12_528  = SUM(( (din_a[151] & din_b[149]) ) + ( Xd_0__inst_mult_12_518  ) + ( Xd_0__inst_mult_12_517  ))
// Xd_0__inst_mult_12_529  = CARRY(( (din_a[151] & din_b[149]) ) + ( Xd_0__inst_mult_12_518  ) + ( Xd_0__inst_mult_12_517  ))
// Xd_0__inst_mult_12_530  = SHARE((din_a[151] & din_b[150]))

	.dataa(!din_a[151]),
	.datab(!din_b[149]),
	.datac(!din_b[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_517 ),
	.sharein(Xd_0__inst_mult_12_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_528 ),
	.cout(Xd_0__inst_mult_12_529 ),
	.shareout(Xd_0__inst_mult_12_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_155 (
// Equation(s):
// Xd_0__inst_mult_12_532  = SUM(( (din_a[147] & din_b[153]) ) + ( Xd_0__inst_mult_12_522  ) + ( Xd_0__inst_mult_12_521  ))
// Xd_0__inst_mult_12_533  = CARRY(( (din_a[147] & din_b[153]) ) + ( Xd_0__inst_mult_12_522  ) + ( Xd_0__inst_mult_12_521  ))
// Xd_0__inst_mult_12_534  = SHARE((din_a[147] & din_b[154]))

	.dataa(!din_a[147]),
	.datab(!din_b[153]),
	.datac(!din_b[154]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_521 ),
	.sharein(Xd_0__inst_mult_12_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_532 ),
	.cout(Xd_0__inst_mult_12_533 ),
	.shareout(Xd_0__inst_mult_12_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_156 (
// Equation(s):
// Xd_0__inst_mult_12_536  = SUM(( (!din_a[149] & (((din_a[148] & din_b[152])))) # (din_a[149] & (!din_b[151] $ (((!din_a[148]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_526  ) + ( Xd_0__inst_mult_12_525  ))
// Xd_0__inst_mult_12_537  = CARRY(( (!din_a[149] & (((din_a[148] & din_b[152])))) # (din_a[149] & (!din_b[151] $ (((!din_a[148]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_526  ) + ( Xd_0__inst_mult_12_525  ))
// Xd_0__inst_mult_12_538  = SHARE((din_a[149] & (din_b[151] & (din_a[148] & din_b[152]))))

	.dataa(!din_a[149]),
	.datab(!din_b[151]),
	.datac(!din_a[148]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_525 ),
	.sharein(Xd_0__inst_mult_12_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_536 ),
	.cout(Xd_0__inst_mult_12_537 ),
	.shareout(Xd_0__inst_mult_12_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_151 (
// Equation(s):
// Xd_0__inst_mult_13_504  = SUM(( (din_a[163] & din_b[161]) ) + ( Xd_0__inst_mult_13_494  ) + ( Xd_0__inst_mult_13_493  ))
// Xd_0__inst_mult_13_505  = CARRY(( (din_a[163] & din_b[161]) ) + ( Xd_0__inst_mult_13_494  ) + ( Xd_0__inst_mult_13_493  ))
// Xd_0__inst_mult_13_506  = SHARE((din_a[163] & din_b[162]))

	.dataa(!din_a[163]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_493 ),
	.sharein(Xd_0__inst_mult_13_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_504 ),
	.cout(Xd_0__inst_mult_13_505 ),
	.shareout(Xd_0__inst_mult_13_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_152 (
// Equation(s):
// Xd_0__inst_mult_13_508  = SUM(( (din_a[159] & din_b[165]) ) + ( Xd_0__inst_mult_13_498  ) + ( Xd_0__inst_mult_13_497  ))
// Xd_0__inst_mult_13_509  = CARRY(( (din_a[159] & din_b[165]) ) + ( Xd_0__inst_mult_13_498  ) + ( Xd_0__inst_mult_13_497  ))
// Xd_0__inst_mult_13_510  = SHARE((din_a[159] & din_b[166]))

	.dataa(!din_a[159]),
	.datab(!din_b[165]),
	.datac(!din_b[166]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_497 ),
	.sharein(Xd_0__inst_mult_13_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_508 ),
	.cout(Xd_0__inst_mult_13_509 ),
	.shareout(Xd_0__inst_mult_13_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_153 (
// Equation(s):
// Xd_0__inst_mult_13_512  = SUM(( (!din_a[161] & (((din_a[160] & din_b[164])))) # (din_a[161] & (!din_b[163] $ (((!din_a[160]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_502  ) + ( Xd_0__inst_mult_13_501  ))
// Xd_0__inst_mult_13_513  = CARRY(( (!din_a[161] & (((din_a[160] & din_b[164])))) # (din_a[161] & (!din_b[163] $ (((!din_a[160]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_502  ) + ( Xd_0__inst_mult_13_501  ))
// Xd_0__inst_mult_13_514  = SHARE((din_a[161] & (din_b[163] & (din_a[160] & din_b[164]))))

	.dataa(!din_a[161]),
	.datab(!din_b[163]),
	.datac(!din_a[160]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_501 ),
	.sharein(Xd_0__inst_mult_13_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_512 ),
	.cout(Xd_0__inst_mult_13_513 ),
	.shareout(Xd_0__inst_mult_13_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_151 (
// Equation(s):
// Xd_0__inst_mult_14_504  = SUM(( (din_a[175] & din_b[173]) ) + ( Xd_0__inst_mult_14_494  ) + ( Xd_0__inst_mult_14_493  ))
// Xd_0__inst_mult_14_505  = CARRY(( (din_a[175] & din_b[173]) ) + ( Xd_0__inst_mult_14_494  ) + ( Xd_0__inst_mult_14_493  ))
// Xd_0__inst_mult_14_506  = SHARE((din_a[175] & din_b[174]))

	.dataa(!din_a[175]),
	.datab(!din_b[173]),
	.datac(!din_b[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_493 ),
	.sharein(Xd_0__inst_mult_14_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_504 ),
	.cout(Xd_0__inst_mult_14_505 ),
	.shareout(Xd_0__inst_mult_14_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_152 (
// Equation(s):
// Xd_0__inst_mult_14_508  = SUM(( (din_a[171] & din_b[177]) ) + ( Xd_0__inst_mult_14_498  ) + ( Xd_0__inst_mult_14_497  ))
// Xd_0__inst_mult_14_509  = CARRY(( (din_a[171] & din_b[177]) ) + ( Xd_0__inst_mult_14_498  ) + ( Xd_0__inst_mult_14_497  ))
// Xd_0__inst_mult_14_510  = SHARE((din_a[171] & din_b[178]))

	.dataa(!din_a[171]),
	.datab(!din_b[177]),
	.datac(!din_b[178]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_497 ),
	.sharein(Xd_0__inst_mult_14_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_508 ),
	.cout(Xd_0__inst_mult_14_509 ),
	.shareout(Xd_0__inst_mult_14_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_153 (
// Equation(s):
// Xd_0__inst_mult_14_512  = SUM(( (!din_a[173] & (((din_a[172] & din_b[176])))) # (din_a[173] & (!din_b[175] $ (((!din_a[172]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_502  ) + ( Xd_0__inst_mult_14_501  ))
// Xd_0__inst_mult_14_513  = CARRY(( (!din_a[173] & (((din_a[172] & din_b[176])))) # (din_a[173] & (!din_b[175] $ (((!din_a[172]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_502  ) + ( Xd_0__inst_mult_14_501  ))
// Xd_0__inst_mult_14_514  = SHARE((din_a[173] & (din_b[175] & (din_a[172] & din_b[176]))))

	.dataa(!din_a[173]),
	.datab(!din_b[175]),
	.datac(!din_a[172]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_501 ),
	.sharein(Xd_0__inst_mult_14_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_512 ),
	.cout(Xd_0__inst_mult_14_513 ),
	.shareout(Xd_0__inst_mult_14_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_158 (
// Equation(s):
// Xd_0__inst_mult_15_532  = SUM(( (din_a[187] & din_b[185]) ) + ( Xd_0__inst_mult_15_522  ) + ( Xd_0__inst_mult_15_521  ))
// Xd_0__inst_mult_15_533  = CARRY(( (din_a[187] & din_b[185]) ) + ( Xd_0__inst_mult_15_522  ) + ( Xd_0__inst_mult_15_521  ))
// Xd_0__inst_mult_15_534  = SHARE((din_a[187] & din_b[186]))

	.dataa(!din_a[187]),
	.datab(!din_b[185]),
	.datac(!din_b[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_521 ),
	.sharein(Xd_0__inst_mult_15_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_532 ),
	.cout(Xd_0__inst_mult_15_533 ),
	.shareout(Xd_0__inst_mult_15_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_159 (
// Equation(s):
// Xd_0__inst_mult_15_536  = SUM(( (din_a[183] & din_b[189]) ) + ( Xd_0__inst_mult_15_526  ) + ( Xd_0__inst_mult_15_525  ))
// Xd_0__inst_mult_15_537  = CARRY(( (din_a[183] & din_b[189]) ) + ( Xd_0__inst_mult_15_526  ) + ( Xd_0__inst_mult_15_525  ))
// Xd_0__inst_mult_15_538  = SHARE((din_a[183] & din_b[190]))

	.dataa(!din_a[183]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_525 ),
	.sharein(Xd_0__inst_mult_15_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_536 ),
	.cout(Xd_0__inst_mult_15_537 ),
	.shareout(Xd_0__inst_mult_15_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_160 (
// Equation(s):
// Xd_0__inst_mult_15_540  = SUM(( (!din_a[185] & (((din_a[184] & din_b[188])))) # (din_a[185] & (!din_b[187] $ (((!din_a[184]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_530  ) + ( Xd_0__inst_mult_15_529  ))
// Xd_0__inst_mult_15_541  = CARRY(( (!din_a[185] & (((din_a[184] & din_b[188])))) # (din_a[185] & (!din_b[187] $ (((!din_a[184]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_530  ) + ( Xd_0__inst_mult_15_529  ))
// Xd_0__inst_mult_15_542  = SHARE((din_a[185] & (din_b[187] & (din_a[184] & din_b[188]))))

	.dataa(!din_a[185]),
	.datab(!din_b[187]),
	.datac(!din_a[184]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_529 ),
	.sharein(Xd_0__inst_mult_15_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_540 ),
	.cout(Xd_0__inst_mult_15_541 ),
	.shareout(Xd_0__inst_mult_15_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_147 (
// Equation(s):
// Xd_0__inst_mult_10_500  = SUM(( (din_a[127] & din_b[125]) ) + ( Xd_0__inst_mult_10_490  ) + ( Xd_0__inst_mult_10_489  ))
// Xd_0__inst_mult_10_501  = CARRY(( (din_a[127] & din_b[125]) ) + ( Xd_0__inst_mult_10_490  ) + ( Xd_0__inst_mult_10_489  ))
// Xd_0__inst_mult_10_502  = SHARE((din_a[127] & din_b[126]))

	.dataa(!din_a[127]),
	.datab(!din_b[125]),
	.datac(!din_b[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_489 ),
	.sharein(Xd_0__inst_mult_10_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_500 ),
	.cout(Xd_0__inst_mult_10_501 ),
	.shareout(Xd_0__inst_mult_10_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_148 (
// Equation(s):
// Xd_0__inst_mult_10_504  = SUM(( (din_a[123] & din_b[129]) ) + ( Xd_0__inst_mult_10_494  ) + ( Xd_0__inst_mult_10_493  ))
// Xd_0__inst_mult_10_505  = CARRY(( (din_a[123] & din_b[129]) ) + ( Xd_0__inst_mult_10_494  ) + ( Xd_0__inst_mult_10_493  ))
// Xd_0__inst_mult_10_506  = SHARE((din_a[123] & din_b[130]))

	.dataa(!din_a[123]),
	.datab(!din_b[129]),
	.datac(!din_b[130]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_493 ),
	.sharein(Xd_0__inst_mult_10_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_504 ),
	.cout(Xd_0__inst_mult_10_505 ),
	.shareout(Xd_0__inst_mult_10_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_149 (
// Equation(s):
// Xd_0__inst_mult_10_508  = SUM(( (!din_a[125] & (((din_a[124] & din_b[128])))) # (din_a[125] & (!din_b[127] $ (((!din_a[124]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_498  ) + ( Xd_0__inst_mult_10_497  ))
// Xd_0__inst_mult_10_509  = CARRY(( (!din_a[125] & (((din_a[124] & din_b[128])))) # (din_a[125] & (!din_b[127] $ (((!din_a[124]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_498  ) + ( Xd_0__inst_mult_10_497  ))
// Xd_0__inst_mult_10_510  = SHARE((din_a[125] & (din_b[127] & (din_a[124] & din_b[128]))))

	.dataa(!din_a[125]),
	.datab(!din_b[127]),
	.datac(!din_a[124]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_497 ),
	.sharein(Xd_0__inst_mult_10_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_508 ),
	.cout(Xd_0__inst_mult_10_509 ),
	.shareout(Xd_0__inst_mult_10_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_151 (
// Equation(s):
// Xd_0__inst_mult_11_504  = SUM(( (din_a[139] & din_b[137]) ) + ( Xd_0__inst_mult_11_494  ) + ( Xd_0__inst_mult_11_493  ))
// Xd_0__inst_mult_11_505  = CARRY(( (din_a[139] & din_b[137]) ) + ( Xd_0__inst_mult_11_494  ) + ( Xd_0__inst_mult_11_493  ))
// Xd_0__inst_mult_11_506  = SHARE((din_a[139] & din_b[138]))

	.dataa(!din_a[139]),
	.datab(!din_b[137]),
	.datac(!din_b[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_493 ),
	.sharein(Xd_0__inst_mult_11_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_504 ),
	.cout(Xd_0__inst_mult_11_505 ),
	.shareout(Xd_0__inst_mult_11_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_152 (
// Equation(s):
// Xd_0__inst_mult_11_508  = SUM(( (din_a[135] & din_b[141]) ) + ( Xd_0__inst_mult_11_498  ) + ( Xd_0__inst_mult_11_497  ))
// Xd_0__inst_mult_11_509  = CARRY(( (din_a[135] & din_b[141]) ) + ( Xd_0__inst_mult_11_498  ) + ( Xd_0__inst_mult_11_497  ))
// Xd_0__inst_mult_11_510  = SHARE((din_a[135] & din_b[142]))

	.dataa(!din_a[135]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_497 ),
	.sharein(Xd_0__inst_mult_11_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_508 ),
	.cout(Xd_0__inst_mult_11_509 ),
	.shareout(Xd_0__inst_mult_11_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_153 (
// Equation(s):
// Xd_0__inst_mult_11_512  = SUM(( (!din_a[137] & (((din_a[136] & din_b[140])))) # (din_a[137] & (!din_b[139] $ (((!din_a[136]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_502  ) + ( Xd_0__inst_mult_11_501  ))
// Xd_0__inst_mult_11_513  = CARRY(( (!din_a[137] & (((din_a[136] & din_b[140])))) # (din_a[137] & (!din_b[139] $ (((!din_a[136]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_502  ) + ( Xd_0__inst_mult_11_501  ))
// Xd_0__inst_mult_11_514  = SHARE((din_a[137] & (din_b[139] & (din_a[136] & din_b[140]))))

	.dataa(!din_a[137]),
	.datab(!din_b[139]),
	.datac(!din_a[136]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_501 ),
	.sharein(Xd_0__inst_mult_11_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_512 ),
	.cout(Xd_0__inst_mult_11_513 ),
	.shareout(Xd_0__inst_mult_11_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_151 (
// Equation(s):
// Xd_0__inst_mult_8_504  = SUM(( (din_a[103] & din_b[101]) ) + ( Xd_0__inst_mult_8_494  ) + ( Xd_0__inst_mult_8_493  ))
// Xd_0__inst_mult_8_505  = CARRY(( (din_a[103] & din_b[101]) ) + ( Xd_0__inst_mult_8_494  ) + ( Xd_0__inst_mult_8_493  ))
// Xd_0__inst_mult_8_506  = SHARE((din_a[103] & din_b[102]))

	.dataa(!din_a[103]),
	.datab(!din_b[101]),
	.datac(!din_b[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_493 ),
	.sharein(Xd_0__inst_mult_8_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_504 ),
	.cout(Xd_0__inst_mult_8_505 ),
	.shareout(Xd_0__inst_mult_8_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_152 (
// Equation(s):
// Xd_0__inst_mult_8_508  = SUM(( (din_a[99] & din_b[105]) ) + ( Xd_0__inst_mult_8_498  ) + ( Xd_0__inst_mult_8_497  ))
// Xd_0__inst_mult_8_509  = CARRY(( (din_a[99] & din_b[105]) ) + ( Xd_0__inst_mult_8_498  ) + ( Xd_0__inst_mult_8_497  ))
// Xd_0__inst_mult_8_510  = SHARE((din_a[99] & din_b[106]))

	.dataa(!din_a[99]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_497 ),
	.sharein(Xd_0__inst_mult_8_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_508 ),
	.cout(Xd_0__inst_mult_8_509 ),
	.shareout(Xd_0__inst_mult_8_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_153 (
// Equation(s):
// Xd_0__inst_mult_8_512  = SUM(( (!din_a[101] & (((din_a[100] & din_b[104])))) # (din_a[101] & (!din_b[103] $ (((!din_a[100]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_502  ) + ( Xd_0__inst_mult_8_501  ))
// Xd_0__inst_mult_8_513  = CARRY(( (!din_a[101] & (((din_a[100] & din_b[104])))) # (din_a[101] & (!din_b[103] $ (((!din_a[100]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_502  ) + ( Xd_0__inst_mult_8_501  ))
// Xd_0__inst_mult_8_514  = SHARE((din_a[101] & (din_b[103] & (din_a[100] & din_b[104]))))

	.dataa(!din_a[101]),
	.datab(!din_b[103]),
	.datac(!din_a[100]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_501 ),
	.sharein(Xd_0__inst_mult_8_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_512 ),
	.cout(Xd_0__inst_mult_8_513 ),
	.shareout(Xd_0__inst_mult_8_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_147 (
// Equation(s):
// Xd_0__inst_mult_9_500  = SUM(( (din_a[115] & din_b[113]) ) + ( Xd_0__inst_mult_9_490  ) + ( Xd_0__inst_mult_9_489  ))
// Xd_0__inst_mult_9_501  = CARRY(( (din_a[115] & din_b[113]) ) + ( Xd_0__inst_mult_9_490  ) + ( Xd_0__inst_mult_9_489  ))
// Xd_0__inst_mult_9_502  = SHARE((din_a[115] & din_b[114]))

	.dataa(!din_a[115]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_489 ),
	.sharein(Xd_0__inst_mult_9_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_500 ),
	.cout(Xd_0__inst_mult_9_501 ),
	.shareout(Xd_0__inst_mult_9_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_148 (
// Equation(s):
// Xd_0__inst_mult_9_504  = SUM(( (din_a[111] & din_b[117]) ) + ( Xd_0__inst_mult_9_494  ) + ( Xd_0__inst_mult_9_493  ))
// Xd_0__inst_mult_9_505  = CARRY(( (din_a[111] & din_b[117]) ) + ( Xd_0__inst_mult_9_494  ) + ( Xd_0__inst_mult_9_493  ))
// Xd_0__inst_mult_9_506  = SHARE((din_a[111] & din_b[118]))

	.dataa(!din_a[111]),
	.datab(!din_b[117]),
	.datac(!din_b[118]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_493 ),
	.sharein(Xd_0__inst_mult_9_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_504 ),
	.cout(Xd_0__inst_mult_9_505 ),
	.shareout(Xd_0__inst_mult_9_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_149 (
// Equation(s):
// Xd_0__inst_mult_9_508  = SUM(( (!din_a[113] & (((din_a[112] & din_b[116])))) # (din_a[113] & (!din_b[115] $ (((!din_a[112]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_498  ) + ( Xd_0__inst_mult_9_497  ))
// Xd_0__inst_mult_9_509  = CARRY(( (!din_a[113] & (((din_a[112] & din_b[116])))) # (din_a[113] & (!din_b[115] $ (((!din_a[112]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_498  ) + ( Xd_0__inst_mult_9_497  ))
// Xd_0__inst_mult_9_510  = SHARE((din_a[113] & (din_b[115] & (din_a[112] & din_b[116]))))

	.dataa(!din_a[113]),
	.datab(!din_b[115]),
	.datac(!din_a[112]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_497 ),
	.sharein(Xd_0__inst_mult_9_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_508 ),
	.cout(Xd_0__inst_mult_9_509 ),
	.shareout(Xd_0__inst_mult_9_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_147 (
// Equation(s):
// Xd_0__inst_mult_6_500  = SUM(( (din_a[79] & din_b[77]) ) + ( Xd_0__inst_mult_6_490  ) + ( Xd_0__inst_mult_6_489  ))
// Xd_0__inst_mult_6_501  = CARRY(( (din_a[79] & din_b[77]) ) + ( Xd_0__inst_mult_6_490  ) + ( Xd_0__inst_mult_6_489  ))
// Xd_0__inst_mult_6_502  = SHARE((din_a[79] & din_b[78]))

	.dataa(!din_a[79]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_489 ),
	.sharein(Xd_0__inst_mult_6_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_500 ),
	.cout(Xd_0__inst_mult_6_501 ),
	.shareout(Xd_0__inst_mult_6_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_148 (
// Equation(s):
// Xd_0__inst_mult_6_504  = SUM(( (din_a[75] & din_b[81]) ) + ( Xd_0__inst_mult_6_494  ) + ( Xd_0__inst_mult_6_493  ))
// Xd_0__inst_mult_6_505  = CARRY(( (din_a[75] & din_b[81]) ) + ( Xd_0__inst_mult_6_494  ) + ( Xd_0__inst_mult_6_493  ))
// Xd_0__inst_mult_6_506  = SHARE((din_a[75] & din_b[82]))

	.dataa(!din_a[75]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_493 ),
	.sharein(Xd_0__inst_mult_6_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_504 ),
	.cout(Xd_0__inst_mult_6_505 ),
	.shareout(Xd_0__inst_mult_6_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_149 (
// Equation(s):
// Xd_0__inst_mult_6_508  = SUM(( (!din_a[77] & (((din_a[76] & din_b[80])))) # (din_a[77] & (!din_b[79] $ (((!din_a[76]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_498  ) + ( Xd_0__inst_mult_6_497  ))
// Xd_0__inst_mult_6_509  = CARRY(( (!din_a[77] & (((din_a[76] & din_b[80])))) # (din_a[77] & (!din_b[79] $ (((!din_a[76]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_498  ) + ( Xd_0__inst_mult_6_497  ))
// Xd_0__inst_mult_6_510  = SHARE((din_a[77] & (din_b[79] & (din_a[76] & din_b[80]))))

	.dataa(!din_a[77]),
	.datab(!din_b[79]),
	.datac(!din_a[76]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_497 ),
	.sharein(Xd_0__inst_mult_6_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_508 ),
	.cout(Xd_0__inst_mult_6_509 ),
	.shareout(Xd_0__inst_mult_6_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_143 (
// Equation(s):
// Xd_0__inst_mult_7_484  = SUM(( GND ) + ( Xd_0__inst_mult_7_466  ) + ( Xd_0__inst_mult_7_465  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_465 ),
	.sharein(Xd_0__inst_mult_7_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_484 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_144 (
// Equation(s):
// Xd_0__inst_mult_7_488  = SUM(( (!din_a[93] & (((din_a[92] & din_b[88])))) # (din_a[93] & (!din_b[87] $ (((!din_a[92]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_470  ) + ( Xd_0__inst_mult_7_469  ))
// Xd_0__inst_mult_7_489  = CARRY(( (!din_a[93] & (((din_a[92] & din_b[88])))) # (din_a[93] & (!din_b[87] $ (((!din_a[92]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_470  ) + ( Xd_0__inst_mult_7_469  ))
// Xd_0__inst_mult_7_490  = SHARE((din_a[93] & (din_b[87] & (din_a[92] & din_b[88]))))

	.dataa(!din_a[93]),
	.datab(!din_b[87]),
	.datac(!din_a[92]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_469 ),
	.sharein(Xd_0__inst_mult_7_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_488 ),
	.cout(Xd_0__inst_mult_7_489 ),
	.shareout(Xd_0__inst_mult_7_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_145 (
// Equation(s):
// Xd_0__inst_mult_7_492  = SUM(( (din_a[91] & din_b[89]) ) + ( Xd_0__inst_mult_7_474  ) + ( Xd_0__inst_mult_7_473  ))
// Xd_0__inst_mult_7_493  = CARRY(( (din_a[91] & din_b[89]) ) + ( Xd_0__inst_mult_7_474  ) + ( Xd_0__inst_mult_7_473  ))
// Xd_0__inst_mult_7_494  = SHARE((din_a[91] & din_b[90]))

	.dataa(!din_a[91]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_473 ),
	.sharein(Xd_0__inst_mult_7_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_492 ),
	.cout(Xd_0__inst_mult_7_493 ),
	.shareout(Xd_0__inst_mult_7_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_146 (
// Equation(s):
// Xd_0__inst_mult_7_496  = SUM(( (din_a[87] & din_b[93]) ) + ( Xd_0__inst_mult_7_478  ) + ( Xd_0__inst_mult_7_477  ))
// Xd_0__inst_mult_7_497  = CARRY(( (din_a[87] & din_b[93]) ) + ( Xd_0__inst_mult_7_478  ) + ( Xd_0__inst_mult_7_477  ))
// Xd_0__inst_mult_7_498  = SHARE((din_a[87] & din_b[94]))

	.dataa(!din_a[87]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_477 ),
	.sharein(Xd_0__inst_mult_7_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_496 ),
	.cout(Xd_0__inst_mult_7_497 ),
	.shareout(Xd_0__inst_mult_7_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_147 (
// Equation(s):
// Xd_0__inst_mult_7_500  = SUM(( (!din_a[89] & (((din_a[88] & din_b[92])))) # (din_a[89] & (!din_b[91] $ (((!din_a[88]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_482  ) + ( Xd_0__inst_mult_7_481  ))
// Xd_0__inst_mult_7_501  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[92])))) # (din_a[89] & (!din_b[91] $ (((!din_a[88]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_482  ) + ( Xd_0__inst_mult_7_481  ))
// Xd_0__inst_mult_7_502  = SHARE((din_a[89] & (din_b[91] & (din_a[88] & din_b[92]))))

	.dataa(!din_a[89]),
	.datab(!din_b[91]),
	.datac(!din_a[88]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_481 ),
	.sharein(Xd_0__inst_mult_7_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_500 ),
	.cout(Xd_0__inst_mult_7_501 ),
	.shareout(Xd_0__inst_mult_7_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_155 (
// Equation(s):
// Xd_0__inst_mult_4_520  = SUM(( GND ) + ( Xd_0__inst_mult_4_506  ) + ( Xd_0__inst_mult_4_505  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_505 ),
	.sharein(Xd_0__inst_mult_4_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_520 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_156 (
// Equation(s):
// Xd_0__inst_mult_4_524  = SUM(( (!din_a[57] & (((din_a[56] & din_b[52])))) # (din_a[57] & (!din_b[51] $ (((!din_a[56]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_510  ) + ( Xd_0__inst_mult_4_509  ))
// Xd_0__inst_mult_4_525  = CARRY(( (!din_a[57] & (((din_a[56] & din_b[52])))) # (din_a[57] & (!din_b[51] $ (((!din_a[56]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_510  ) + ( Xd_0__inst_mult_4_509  ))
// Xd_0__inst_mult_4_526  = SHARE((din_a[57] & (din_b[51] & (din_a[56] & din_b[52]))))

	.dataa(!din_a[57]),
	.datab(!din_b[51]),
	.datac(!din_a[56]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_509 ),
	.sharein(Xd_0__inst_mult_4_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_524 ),
	.cout(Xd_0__inst_mult_4_525 ),
	.shareout(Xd_0__inst_mult_4_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_157 (
// Equation(s):
// Xd_0__inst_mult_4_528  = SUM(( (din_a[55] & din_b[53]) ) + ( Xd_0__inst_mult_4_514  ) + ( Xd_0__inst_mult_4_513  ))
// Xd_0__inst_mult_4_529  = CARRY(( (din_a[55] & din_b[53]) ) + ( Xd_0__inst_mult_4_514  ) + ( Xd_0__inst_mult_4_513  ))
// Xd_0__inst_mult_4_530  = SHARE((din_a[55] & din_b[54]))

	.dataa(!din_a[55]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_513 ),
	.sharein(Xd_0__inst_mult_4_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_528 ),
	.cout(Xd_0__inst_mult_4_529 ),
	.shareout(Xd_0__inst_mult_4_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_158 (
// Equation(s):
// Xd_0__inst_mult_4_532  = SUM(( (!din_a[53] & (((din_a[52] & din_b[56])))) # (din_a[53] & (!din_b[55] $ (((!din_a[52]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_518  ) + ( Xd_0__inst_mult_4_517  ))
// Xd_0__inst_mult_4_533  = CARRY(( (!din_a[53] & (((din_a[52] & din_b[56])))) # (din_a[53] & (!din_b[55] $ (((!din_a[52]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_518  ) + ( Xd_0__inst_mult_4_517  ))
// Xd_0__inst_mult_4_534  = SHARE((din_a[53] & (din_b[55] & (din_a[52] & din_b[56]))))

	.dataa(!din_a[53]),
	.datab(!din_b[55]),
	.datac(!din_a[52]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_517 ),
	.sharein(Xd_0__inst_mult_4_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_532 ),
	.cout(Xd_0__inst_mult_4_533 ),
	.shareout(Xd_0__inst_mult_4_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_143 (
// Equation(s):
// Xd_0__inst_mult_5_484  = SUM(( GND ) + ( Xd_0__inst_mult_5_466  ) + ( Xd_0__inst_mult_5_465  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_465 ),
	.sharein(Xd_0__inst_mult_5_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_484 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_144 (
// Equation(s):
// Xd_0__inst_mult_5_488  = SUM(( (!din_a[69] & (((din_a[68] & din_b[64])))) # (din_a[69] & (!din_b[63] $ (((!din_a[68]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_470  ) + ( Xd_0__inst_mult_5_469  ))
// Xd_0__inst_mult_5_489  = CARRY(( (!din_a[69] & (((din_a[68] & din_b[64])))) # (din_a[69] & (!din_b[63] $ (((!din_a[68]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_470  ) + ( Xd_0__inst_mult_5_469  ))
// Xd_0__inst_mult_5_490  = SHARE((din_a[69] & (din_b[63] & (din_a[68] & din_b[64]))))

	.dataa(!din_a[69]),
	.datab(!din_b[63]),
	.datac(!din_a[68]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_469 ),
	.sharein(Xd_0__inst_mult_5_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_488 ),
	.cout(Xd_0__inst_mult_5_489 ),
	.shareout(Xd_0__inst_mult_5_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_145 (
// Equation(s):
// Xd_0__inst_mult_5_492  = SUM(( (din_a[67] & din_b[65]) ) + ( Xd_0__inst_mult_5_474  ) + ( Xd_0__inst_mult_5_473  ))
// Xd_0__inst_mult_5_493  = CARRY(( (din_a[67] & din_b[65]) ) + ( Xd_0__inst_mult_5_474  ) + ( Xd_0__inst_mult_5_473  ))
// Xd_0__inst_mult_5_494  = SHARE((din_a[67] & din_b[66]))

	.dataa(!din_a[67]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_473 ),
	.sharein(Xd_0__inst_mult_5_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_492 ),
	.cout(Xd_0__inst_mult_5_493 ),
	.shareout(Xd_0__inst_mult_5_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_146 (
// Equation(s):
// Xd_0__inst_mult_5_496  = SUM(( (din_a[63] & din_b[69]) ) + ( Xd_0__inst_mult_5_478  ) + ( Xd_0__inst_mult_5_477  ))
// Xd_0__inst_mult_5_497  = CARRY(( (din_a[63] & din_b[69]) ) + ( Xd_0__inst_mult_5_478  ) + ( Xd_0__inst_mult_5_477  ))
// Xd_0__inst_mult_5_498  = SHARE((din_a[63] & din_b[70]))

	.dataa(!din_a[63]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_477 ),
	.sharein(Xd_0__inst_mult_5_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_496 ),
	.cout(Xd_0__inst_mult_5_497 ),
	.shareout(Xd_0__inst_mult_5_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_147 (
// Equation(s):
// Xd_0__inst_mult_5_500  = SUM(( (!din_a[65] & (((din_a[64] & din_b[68])))) # (din_a[65] & (!din_b[67] $ (((!din_a[64]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_482  ) + ( Xd_0__inst_mult_5_481  ))
// Xd_0__inst_mult_5_501  = CARRY(( (!din_a[65] & (((din_a[64] & din_b[68])))) # (din_a[65] & (!din_b[67] $ (((!din_a[64]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_482  ) + ( Xd_0__inst_mult_5_481  ))
// Xd_0__inst_mult_5_502  = SHARE((din_a[65] & (din_b[67] & (din_a[64] & din_b[68]))))

	.dataa(!din_a[65]),
	.datab(!din_b[67]),
	.datac(!din_a[64]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_481 ),
	.sharein(Xd_0__inst_mult_5_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_500 ),
	.cout(Xd_0__inst_mult_5_501 ),
	.shareout(Xd_0__inst_mult_5_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_147 (
// Equation(s):
// Xd_0__inst_mult_2_488  = SUM(( GND ) + ( Xd_0__inst_mult_2_470  ) + ( Xd_0__inst_mult_2_469  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_469 ),
	.sharein(Xd_0__inst_mult_2_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_488 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_148 (
// Equation(s):
// Xd_0__inst_mult_2_492  = SUM(( (!din_a[33] & (((din_a[32] & din_b[28])))) # (din_a[33] & (!din_b[27] $ (((!din_a[32]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_474  ) + ( Xd_0__inst_mult_2_473  ))
// Xd_0__inst_mult_2_493  = CARRY(( (!din_a[33] & (((din_a[32] & din_b[28])))) # (din_a[33] & (!din_b[27] $ (((!din_a[32]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_474  ) + ( Xd_0__inst_mult_2_473  ))
// Xd_0__inst_mult_2_494  = SHARE((din_a[33] & (din_b[27] & (din_a[32] & din_b[28]))))

	.dataa(!din_a[33]),
	.datab(!din_b[27]),
	.datac(!din_a[32]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_473 ),
	.sharein(Xd_0__inst_mult_2_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_492 ),
	.cout(Xd_0__inst_mult_2_493 ),
	.shareout(Xd_0__inst_mult_2_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_149 (
// Equation(s):
// Xd_0__inst_mult_2_496  = SUM(( (din_a[31] & din_b[29]) ) + ( Xd_0__inst_mult_2_478  ) + ( Xd_0__inst_mult_2_477  ))
// Xd_0__inst_mult_2_497  = CARRY(( (din_a[31] & din_b[29]) ) + ( Xd_0__inst_mult_2_478  ) + ( Xd_0__inst_mult_2_477  ))
// Xd_0__inst_mult_2_498  = SHARE((din_a[31] & din_b[30]))

	.dataa(!din_a[31]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_477 ),
	.sharein(Xd_0__inst_mult_2_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_496 ),
	.cout(Xd_0__inst_mult_2_497 ),
	.shareout(Xd_0__inst_mult_2_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_150 (
// Equation(s):
// Xd_0__inst_mult_2_500  = SUM(( (din_a[27] & din_b[33]) ) + ( Xd_0__inst_mult_2_482  ) + ( Xd_0__inst_mult_2_481  ))
// Xd_0__inst_mult_2_501  = CARRY(( (din_a[27] & din_b[33]) ) + ( Xd_0__inst_mult_2_482  ) + ( Xd_0__inst_mult_2_481  ))
// Xd_0__inst_mult_2_502  = SHARE((din_a[27] & din_b[34]))

	.dataa(!din_a[27]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_481 ),
	.sharein(Xd_0__inst_mult_2_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_500 ),
	.cout(Xd_0__inst_mult_2_501 ),
	.shareout(Xd_0__inst_mult_2_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_151 (
// Equation(s):
// Xd_0__inst_mult_2_504  = SUM(( (!din_a[29] & (((din_a[28] & din_b[32])))) # (din_a[29] & (!din_b[31] $ (((!din_a[28]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_486  ) + ( Xd_0__inst_mult_2_485  ))
// Xd_0__inst_mult_2_505  = CARRY(( (!din_a[29] & (((din_a[28] & din_b[32])))) # (din_a[29] & (!din_b[31] $ (((!din_a[28]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_486  ) + ( Xd_0__inst_mult_2_485  ))
// Xd_0__inst_mult_2_506  = SHARE((din_a[29] & (din_b[31] & (din_a[28] & din_b[32]))))

	.dataa(!din_a[29]),
	.datab(!din_b[31]),
	.datac(!din_a[28]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_485 ),
	.sharein(Xd_0__inst_mult_2_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_504 ),
	.cout(Xd_0__inst_mult_2_505 ),
	.shareout(Xd_0__inst_mult_2_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_143 (
// Equation(s):
// Xd_0__inst_mult_3_484  = SUM(( GND ) + ( Xd_0__inst_mult_3_466  ) + ( Xd_0__inst_mult_3_465  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_465 ),
	.sharein(Xd_0__inst_mult_3_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_484 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_144 (
// Equation(s):
// Xd_0__inst_mult_3_488  = SUM(( (!din_a[45] & (((din_a[44] & din_b[40])))) # (din_a[45] & (!din_b[39] $ (((!din_a[44]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_470  ) + ( Xd_0__inst_mult_3_469  ))
// Xd_0__inst_mult_3_489  = CARRY(( (!din_a[45] & (((din_a[44] & din_b[40])))) # (din_a[45] & (!din_b[39] $ (((!din_a[44]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_470  ) + ( Xd_0__inst_mult_3_469  ))
// Xd_0__inst_mult_3_490  = SHARE((din_a[45] & (din_b[39] & (din_a[44] & din_b[40]))))

	.dataa(!din_a[45]),
	.datab(!din_b[39]),
	.datac(!din_a[44]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_469 ),
	.sharein(Xd_0__inst_mult_3_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_488 ),
	.cout(Xd_0__inst_mult_3_489 ),
	.shareout(Xd_0__inst_mult_3_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_145 (
// Equation(s):
// Xd_0__inst_mult_3_492  = SUM(( (din_a[43] & din_b[41]) ) + ( Xd_0__inst_mult_3_474  ) + ( Xd_0__inst_mult_3_473  ))
// Xd_0__inst_mult_3_493  = CARRY(( (din_a[43] & din_b[41]) ) + ( Xd_0__inst_mult_3_474  ) + ( Xd_0__inst_mult_3_473  ))
// Xd_0__inst_mult_3_494  = SHARE((din_a[43] & din_b[42]))

	.dataa(!din_a[43]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_473 ),
	.sharein(Xd_0__inst_mult_3_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_492 ),
	.cout(Xd_0__inst_mult_3_493 ),
	.shareout(Xd_0__inst_mult_3_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_146 (
// Equation(s):
// Xd_0__inst_mult_3_496  = SUM(( (din_a[39] & din_b[45]) ) + ( Xd_0__inst_mult_3_478  ) + ( Xd_0__inst_mult_3_477  ))
// Xd_0__inst_mult_3_497  = CARRY(( (din_a[39] & din_b[45]) ) + ( Xd_0__inst_mult_3_478  ) + ( Xd_0__inst_mult_3_477  ))
// Xd_0__inst_mult_3_498  = SHARE((din_a[39] & din_b[46]))

	.dataa(!din_a[39]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_477 ),
	.sharein(Xd_0__inst_mult_3_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_496 ),
	.cout(Xd_0__inst_mult_3_497 ),
	.shareout(Xd_0__inst_mult_3_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_147 (
// Equation(s):
// Xd_0__inst_mult_3_500  = SUM(( (!din_a[41] & (((din_a[40] & din_b[44])))) # (din_a[41] & (!din_b[43] $ (((!din_a[40]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_482  ) + ( Xd_0__inst_mult_3_481  ))
// Xd_0__inst_mult_3_501  = CARRY(( (!din_a[41] & (((din_a[40] & din_b[44])))) # (din_a[41] & (!din_b[43] $ (((!din_a[40]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_482  ) + ( Xd_0__inst_mult_3_481  ))
// Xd_0__inst_mult_3_502  = SHARE((din_a[41] & (din_b[43] & (din_a[40] & din_b[44]))))

	.dataa(!din_a[41]),
	.datab(!din_b[43]),
	.datac(!din_a[40]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_481 ),
	.sharein(Xd_0__inst_mult_3_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_500 ),
	.cout(Xd_0__inst_mult_3_501 ),
	.shareout(Xd_0__inst_mult_3_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_147 (
// Equation(s):
// Xd_0__inst_mult_0_488  = SUM(( GND ) + ( Xd_0__inst_mult_0_470  ) + ( Xd_0__inst_mult_0_469  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_469 ),
	.sharein(Xd_0__inst_mult_0_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_488 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_148 (
// Equation(s):
// Xd_0__inst_mult_0_492  = SUM(( (!din_a[9] & (((din_a[8] & din_b[4])))) # (din_a[9] & (!din_b[3] $ (((!din_a[8]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_474  ) + ( Xd_0__inst_mult_0_473  ))
// Xd_0__inst_mult_0_493  = CARRY(( (!din_a[9] & (((din_a[8] & din_b[4])))) # (din_a[9] & (!din_b[3] $ (((!din_a[8]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_474  ) + ( Xd_0__inst_mult_0_473  ))
// Xd_0__inst_mult_0_494  = SHARE((din_a[9] & (din_b[3] & (din_a[8] & din_b[4]))))

	.dataa(!din_a[9]),
	.datab(!din_b[3]),
	.datac(!din_a[8]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_473 ),
	.sharein(Xd_0__inst_mult_0_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_492 ),
	.cout(Xd_0__inst_mult_0_493 ),
	.shareout(Xd_0__inst_mult_0_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_149 (
// Equation(s):
// Xd_0__inst_mult_0_496  = SUM(( (din_a[7] & din_b[5]) ) + ( Xd_0__inst_mult_0_478  ) + ( Xd_0__inst_mult_0_477  ))
// Xd_0__inst_mult_0_497  = CARRY(( (din_a[7] & din_b[5]) ) + ( Xd_0__inst_mult_0_478  ) + ( Xd_0__inst_mult_0_477  ))
// Xd_0__inst_mult_0_498  = SHARE((din_a[7] & din_b[6]))

	.dataa(!din_a[7]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_477 ),
	.sharein(Xd_0__inst_mult_0_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_496 ),
	.cout(Xd_0__inst_mult_0_497 ),
	.shareout(Xd_0__inst_mult_0_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_150 (
// Equation(s):
// Xd_0__inst_mult_0_500  = SUM(( (din_a[3] & din_b[9]) ) + ( Xd_0__inst_mult_0_482  ) + ( Xd_0__inst_mult_0_481  ))
// Xd_0__inst_mult_0_501  = CARRY(( (din_a[3] & din_b[9]) ) + ( Xd_0__inst_mult_0_482  ) + ( Xd_0__inst_mult_0_481  ))
// Xd_0__inst_mult_0_502  = SHARE((din_a[3] & din_b[10]))

	.dataa(!din_a[3]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_481 ),
	.sharein(Xd_0__inst_mult_0_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_500 ),
	.cout(Xd_0__inst_mult_0_501 ),
	.shareout(Xd_0__inst_mult_0_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_151 (
// Equation(s):
// Xd_0__inst_mult_0_504  = SUM(( (!din_a[5] & (((din_a[4] & din_b[8])))) # (din_a[5] & (!din_b[7] $ (((!din_a[4]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_486  ) + ( Xd_0__inst_mult_0_485  ))
// Xd_0__inst_mult_0_505  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[8])))) # (din_a[5] & (!din_b[7] $ (((!din_a[4]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_486  ) + ( Xd_0__inst_mult_0_485  ))
// Xd_0__inst_mult_0_506  = SHARE((din_a[5] & (din_b[7] & (din_a[4] & din_b[8]))))

	.dataa(!din_a[5]),
	.datab(!din_b[7]),
	.datac(!din_a[4]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_485 ),
	.sharein(Xd_0__inst_mult_0_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_504 ),
	.cout(Xd_0__inst_mult_0_505 ),
	.shareout(Xd_0__inst_mult_0_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_147 (
// Equation(s):
// Xd_0__inst_mult_1_488  = SUM(( GND ) + ( Xd_0__inst_mult_1_470  ) + ( Xd_0__inst_mult_1_469  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_469 ),
	.sharein(Xd_0__inst_mult_1_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_488 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_148 (
// Equation(s):
// Xd_0__inst_mult_1_492  = SUM(( (!din_a[21] & (((din_a[20] & din_b[16])))) # (din_a[21] & (!din_b[15] $ (((!din_a[20]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_474  ) + ( Xd_0__inst_mult_1_473  ))
// Xd_0__inst_mult_1_493  = CARRY(( (!din_a[21] & (((din_a[20] & din_b[16])))) # (din_a[21] & (!din_b[15] $ (((!din_a[20]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_474  ) + ( Xd_0__inst_mult_1_473  ))
// Xd_0__inst_mult_1_494  = SHARE((din_a[21] & (din_b[15] & (din_a[20] & din_b[16]))))

	.dataa(!din_a[21]),
	.datab(!din_b[15]),
	.datac(!din_a[20]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_473 ),
	.sharein(Xd_0__inst_mult_1_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_492 ),
	.cout(Xd_0__inst_mult_1_493 ),
	.shareout(Xd_0__inst_mult_1_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_149 (
// Equation(s):
// Xd_0__inst_mult_1_496  = SUM(( (din_a[19] & din_b[17]) ) + ( Xd_0__inst_mult_1_478  ) + ( Xd_0__inst_mult_1_477  ))
// Xd_0__inst_mult_1_497  = CARRY(( (din_a[19] & din_b[17]) ) + ( Xd_0__inst_mult_1_478  ) + ( Xd_0__inst_mult_1_477  ))
// Xd_0__inst_mult_1_498  = SHARE((din_a[19] & din_b[18]))

	.dataa(!din_a[19]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_477 ),
	.sharein(Xd_0__inst_mult_1_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_496 ),
	.cout(Xd_0__inst_mult_1_497 ),
	.shareout(Xd_0__inst_mult_1_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_150 (
// Equation(s):
// Xd_0__inst_mult_1_500  = SUM(( (din_a[15] & din_b[21]) ) + ( Xd_0__inst_mult_1_482  ) + ( Xd_0__inst_mult_1_481  ))
// Xd_0__inst_mult_1_501  = CARRY(( (din_a[15] & din_b[21]) ) + ( Xd_0__inst_mult_1_482  ) + ( Xd_0__inst_mult_1_481  ))
// Xd_0__inst_mult_1_502  = SHARE((din_a[15] & din_b[22]))

	.dataa(!din_a[15]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_481 ),
	.sharein(Xd_0__inst_mult_1_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_500 ),
	.cout(Xd_0__inst_mult_1_501 ),
	.shareout(Xd_0__inst_mult_1_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_151 (
// Equation(s):
// Xd_0__inst_mult_1_504  = SUM(( (!din_a[17] & (((din_a[16] & din_b[20])))) # (din_a[17] & (!din_b[19] $ (((!din_a[16]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_486  ) + ( Xd_0__inst_mult_1_485  ))
// Xd_0__inst_mult_1_505  = CARRY(( (!din_a[17] & (((din_a[16] & din_b[20])))) # (din_a[17] & (!din_b[19] $ (((!din_a[16]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_486  ) + ( Xd_0__inst_mult_1_485  ))
// Xd_0__inst_mult_1_506  = SHARE((din_a[17] & (din_b[19] & (din_a[16] & din_b[20]))))

	.dataa(!din_a[17]),
	.datab(!din_b[19]),
	.datac(!din_a[16]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_485 ),
	.sharein(Xd_0__inst_mult_1_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_504 ),
	.cout(Xd_0__inst_mult_1_505 ),
	.shareout(Xd_0__inst_mult_1_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_157 (
// Equation(s):
// Xd_0__inst_mult_12_540  = SUM(( (din_a[152] & din_b[149]) ) + ( Xd_0__inst_mult_12_530  ) + ( Xd_0__inst_mult_12_529  ))
// Xd_0__inst_mult_12_541  = CARRY(( (din_a[152] & din_b[149]) ) + ( Xd_0__inst_mult_12_530  ) + ( Xd_0__inst_mult_12_529  ))
// Xd_0__inst_mult_12_542  = SHARE((din_a[152] & din_b[150]))

	.dataa(!din_a[152]),
	.datab(!din_b[149]),
	.datac(!din_b[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_529 ),
	.sharein(Xd_0__inst_mult_12_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_540 ),
	.cout(Xd_0__inst_mult_12_541 ),
	.shareout(Xd_0__inst_mult_12_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_158 (
// Equation(s):
// Xd_0__inst_mult_12_544  = SUM(( (!din_a[150] & (((din_a[149] & din_b[152])))) # (din_a[150] & (!din_b[151] $ (((!din_a[149]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_538  ) + ( Xd_0__inst_mult_12_537  ))
// Xd_0__inst_mult_12_545  = CARRY(( (!din_a[150] & (((din_a[149] & din_b[152])))) # (din_a[150] & (!din_b[151] $ (((!din_a[149]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_538  ) + ( Xd_0__inst_mult_12_537  ))
// Xd_0__inst_mult_12_546  = SHARE((din_a[150] & (din_b[151] & (din_a[149] & din_b[152]))))

	.dataa(!din_a[150]),
	.datab(!din_b[151]),
	.datac(!din_a[149]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_537 ),
	.sharein(Xd_0__inst_mult_12_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_544 ),
	.cout(Xd_0__inst_mult_12_545 ),
	.shareout(Xd_0__inst_mult_12_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_154 (
// Equation(s):
// Xd_0__inst_mult_13_516  = SUM(( (din_a[164] & din_b[161]) ) + ( Xd_0__inst_mult_13_506  ) + ( Xd_0__inst_mult_13_505  ))
// Xd_0__inst_mult_13_517  = CARRY(( (din_a[164] & din_b[161]) ) + ( Xd_0__inst_mult_13_506  ) + ( Xd_0__inst_mult_13_505  ))
// Xd_0__inst_mult_13_518  = SHARE((din_a[164] & din_b[162]))

	.dataa(!din_a[164]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_505 ),
	.sharein(Xd_0__inst_mult_13_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_516 ),
	.cout(Xd_0__inst_mult_13_517 ),
	.shareout(Xd_0__inst_mult_13_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_155 (
// Equation(s):
// Xd_0__inst_mult_13_520  = SUM(( (din_a[160] & din_b[165]) ) + ( Xd_0__inst_mult_13_510  ) + ( Xd_0__inst_mult_13_509  ))
// Xd_0__inst_mult_13_521  = CARRY(( (din_a[160] & din_b[165]) ) + ( Xd_0__inst_mult_13_510  ) + ( Xd_0__inst_mult_13_509  ))
// Xd_0__inst_mult_13_522  = SHARE((din_a[160] & din_b[166]))

	.dataa(!din_a[160]),
	.datab(!din_b[165]),
	.datac(!din_b[166]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_509 ),
	.sharein(Xd_0__inst_mult_13_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_520 ),
	.cout(Xd_0__inst_mult_13_521 ),
	.shareout(Xd_0__inst_mult_13_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_156 (
// Equation(s):
// Xd_0__inst_mult_13_524  = SUM(( (!din_a[162] & (((din_a[161] & din_b[164])))) # (din_a[162] & (!din_b[163] $ (((!din_a[161]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_514  ) + ( Xd_0__inst_mult_13_513  ))
// Xd_0__inst_mult_13_525  = CARRY(( (!din_a[162] & (((din_a[161] & din_b[164])))) # (din_a[162] & (!din_b[163] $ (((!din_a[161]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_514  ) + ( Xd_0__inst_mult_13_513  ))
// Xd_0__inst_mult_13_526  = SHARE((din_a[162] & (din_b[163] & (din_a[161] & din_b[164]))))

	.dataa(!din_a[162]),
	.datab(!din_b[163]),
	.datac(!din_a[161]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_513 ),
	.sharein(Xd_0__inst_mult_13_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_524 ),
	.cout(Xd_0__inst_mult_13_525 ),
	.shareout(Xd_0__inst_mult_13_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_154 (
// Equation(s):
// Xd_0__inst_mult_14_516  = SUM(( (din_a[176] & din_b[173]) ) + ( Xd_0__inst_mult_14_506  ) + ( Xd_0__inst_mult_14_505  ))
// Xd_0__inst_mult_14_517  = CARRY(( (din_a[176] & din_b[173]) ) + ( Xd_0__inst_mult_14_506  ) + ( Xd_0__inst_mult_14_505  ))
// Xd_0__inst_mult_14_518  = SHARE((din_a[176] & din_b[174]))

	.dataa(!din_a[176]),
	.datab(!din_b[173]),
	.datac(!din_b[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_505 ),
	.sharein(Xd_0__inst_mult_14_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_516 ),
	.cout(Xd_0__inst_mult_14_517 ),
	.shareout(Xd_0__inst_mult_14_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_155 (
// Equation(s):
// Xd_0__inst_mult_14_520  = SUM(( (din_a[172] & din_b[177]) ) + ( Xd_0__inst_mult_14_510  ) + ( Xd_0__inst_mult_14_509  ))
// Xd_0__inst_mult_14_521  = CARRY(( (din_a[172] & din_b[177]) ) + ( Xd_0__inst_mult_14_510  ) + ( Xd_0__inst_mult_14_509  ))
// Xd_0__inst_mult_14_522  = SHARE((din_a[172] & din_b[178]))

	.dataa(!din_a[172]),
	.datab(!din_b[177]),
	.datac(!din_b[178]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_509 ),
	.sharein(Xd_0__inst_mult_14_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_520 ),
	.cout(Xd_0__inst_mult_14_521 ),
	.shareout(Xd_0__inst_mult_14_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_156 (
// Equation(s):
// Xd_0__inst_mult_14_524  = SUM(( (!din_a[174] & (((din_a[173] & din_b[176])))) # (din_a[174] & (!din_b[175] $ (((!din_a[173]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_514  ) + ( Xd_0__inst_mult_14_513  ))
// Xd_0__inst_mult_14_525  = CARRY(( (!din_a[174] & (((din_a[173] & din_b[176])))) # (din_a[174] & (!din_b[175] $ (((!din_a[173]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_514  ) + ( Xd_0__inst_mult_14_513  ))
// Xd_0__inst_mult_14_526  = SHARE((din_a[174] & (din_b[175] & (din_a[173] & din_b[176]))))

	.dataa(!din_a[174]),
	.datab(!din_b[175]),
	.datac(!din_a[173]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_513 ),
	.sharein(Xd_0__inst_mult_14_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_524 ),
	.cout(Xd_0__inst_mult_14_525 ),
	.shareout(Xd_0__inst_mult_14_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_161 (
// Equation(s):
// Xd_0__inst_mult_15_544  = SUM(( (din_a[188] & din_b[185]) ) + ( Xd_0__inst_mult_15_534  ) + ( Xd_0__inst_mult_15_533  ))
// Xd_0__inst_mult_15_545  = CARRY(( (din_a[188] & din_b[185]) ) + ( Xd_0__inst_mult_15_534  ) + ( Xd_0__inst_mult_15_533  ))
// Xd_0__inst_mult_15_546  = SHARE((din_a[188] & din_b[186]))

	.dataa(!din_a[188]),
	.datab(!din_b[185]),
	.datac(!din_b[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_533 ),
	.sharein(Xd_0__inst_mult_15_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_544 ),
	.cout(Xd_0__inst_mult_15_545 ),
	.shareout(Xd_0__inst_mult_15_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_162 (
// Equation(s):
// Xd_0__inst_mult_15_548  = SUM(( (!din_a[186] & (((din_a[185] & din_b[188])))) # (din_a[186] & (!din_b[187] $ (((!din_a[185]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_542  ) + ( Xd_0__inst_mult_15_541  ))
// Xd_0__inst_mult_15_549  = CARRY(( (!din_a[186] & (((din_a[185] & din_b[188])))) # (din_a[186] & (!din_b[187] $ (((!din_a[185]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_542  ) + ( Xd_0__inst_mult_15_541  ))
// Xd_0__inst_mult_15_550  = SHARE((din_a[186] & (din_b[187] & (din_a[185] & din_b[188]))))

	.dataa(!din_a[186]),
	.datab(!din_b[187]),
	.datac(!din_a[185]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_541 ),
	.sharein(Xd_0__inst_mult_15_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_548 ),
	.cout(Xd_0__inst_mult_15_549 ),
	.shareout(Xd_0__inst_mult_15_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_150 (
// Equation(s):
// Xd_0__inst_mult_10_512  = SUM(( (din_a[128] & din_b[125]) ) + ( Xd_0__inst_mult_10_502  ) + ( Xd_0__inst_mult_10_501  ))
// Xd_0__inst_mult_10_513  = CARRY(( (din_a[128] & din_b[125]) ) + ( Xd_0__inst_mult_10_502  ) + ( Xd_0__inst_mult_10_501  ))
// Xd_0__inst_mult_10_514  = SHARE((din_a[128] & din_b[126]))

	.dataa(!din_a[128]),
	.datab(!din_b[125]),
	.datac(!din_b[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_501 ),
	.sharein(Xd_0__inst_mult_10_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_512 ),
	.cout(Xd_0__inst_mult_10_513 ),
	.shareout(Xd_0__inst_mult_10_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_151 (
// Equation(s):
// Xd_0__inst_mult_10_516  = SUM(( (din_a[124] & din_b[129]) ) + ( Xd_0__inst_mult_10_506  ) + ( Xd_0__inst_mult_10_505  ))
// Xd_0__inst_mult_10_517  = CARRY(( (din_a[124] & din_b[129]) ) + ( Xd_0__inst_mult_10_506  ) + ( Xd_0__inst_mult_10_505  ))
// Xd_0__inst_mult_10_518  = SHARE((din_a[124] & din_b[130]))

	.dataa(!din_a[124]),
	.datab(!din_b[129]),
	.datac(!din_b[130]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_505 ),
	.sharein(Xd_0__inst_mult_10_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_516 ),
	.cout(Xd_0__inst_mult_10_517 ),
	.shareout(Xd_0__inst_mult_10_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_152 (
// Equation(s):
// Xd_0__inst_mult_10_520  = SUM(( (!din_a[126] & (((din_a[125] & din_b[128])))) # (din_a[126] & (!din_b[127] $ (((!din_a[125]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_510  ) + ( Xd_0__inst_mult_10_509  ))
// Xd_0__inst_mult_10_521  = CARRY(( (!din_a[126] & (((din_a[125] & din_b[128])))) # (din_a[126] & (!din_b[127] $ (((!din_a[125]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_510  ) + ( Xd_0__inst_mult_10_509  ))
// Xd_0__inst_mult_10_522  = SHARE((din_a[126] & (din_b[127] & (din_a[125] & din_b[128]))))

	.dataa(!din_a[126]),
	.datab(!din_b[127]),
	.datac(!din_a[125]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_509 ),
	.sharein(Xd_0__inst_mult_10_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_520 ),
	.cout(Xd_0__inst_mult_10_521 ),
	.shareout(Xd_0__inst_mult_10_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_154 (
// Equation(s):
// Xd_0__inst_mult_11_516  = SUM(( (din_a[140] & din_b[137]) ) + ( Xd_0__inst_mult_11_506  ) + ( Xd_0__inst_mult_11_505  ))
// Xd_0__inst_mult_11_517  = CARRY(( (din_a[140] & din_b[137]) ) + ( Xd_0__inst_mult_11_506  ) + ( Xd_0__inst_mult_11_505  ))
// Xd_0__inst_mult_11_518  = SHARE((din_a[140] & din_b[138]))

	.dataa(!din_a[140]),
	.datab(!din_b[137]),
	.datac(!din_b[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_505 ),
	.sharein(Xd_0__inst_mult_11_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_516 ),
	.cout(Xd_0__inst_mult_11_517 ),
	.shareout(Xd_0__inst_mult_11_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_155 (
// Equation(s):
// Xd_0__inst_mult_11_520  = SUM(( (din_a[136] & din_b[141]) ) + ( Xd_0__inst_mult_11_510  ) + ( Xd_0__inst_mult_11_509  ))
// Xd_0__inst_mult_11_521  = CARRY(( (din_a[136] & din_b[141]) ) + ( Xd_0__inst_mult_11_510  ) + ( Xd_0__inst_mult_11_509  ))
// Xd_0__inst_mult_11_522  = SHARE((din_a[136] & din_b[142]))

	.dataa(!din_a[136]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_509 ),
	.sharein(Xd_0__inst_mult_11_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_520 ),
	.cout(Xd_0__inst_mult_11_521 ),
	.shareout(Xd_0__inst_mult_11_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_156 (
// Equation(s):
// Xd_0__inst_mult_11_524  = SUM(( (!din_a[138] & (((din_a[137] & din_b[140])))) # (din_a[138] & (!din_b[139] $ (((!din_a[137]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_514  ) + ( Xd_0__inst_mult_11_513  ))
// Xd_0__inst_mult_11_525  = CARRY(( (!din_a[138] & (((din_a[137] & din_b[140])))) # (din_a[138] & (!din_b[139] $ (((!din_a[137]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_514  ) + ( Xd_0__inst_mult_11_513  ))
// Xd_0__inst_mult_11_526  = SHARE((din_a[138] & (din_b[139] & (din_a[137] & din_b[140]))))

	.dataa(!din_a[138]),
	.datab(!din_b[139]),
	.datac(!din_a[137]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_513 ),
	.sharein(Xd_0__inst_mult_11_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_524 ),
	.cout(Xd_0__inst_mult_11_525 ),
	.shareout(Xd_0__inst_mult_11_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_154 (
// Equation(s):
// Xd_0__inst_mult_8_516  = SUM(( (din_a[104] & din_b[101]) ) + ( Xd_0__inst_mult_8_506  ) + ( Xd_0__inst_mult_8_505  ))
// Xd_0__inst_mult_8_517  = CARRY(( (din_a[104] & din_b[101]) ) + ( Xd_0__inst_mult_8_506  ) + ( Xd_0__inst_mult_8_505  ))
// Xd_0__inst_mult_8_518  = SHARE((din_a[104] & din_b[102]))

	.dataa(!din_a[104]),
	.datab(!din_b[101]),
	.datac(!din_b[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_505 ),
	.sharein(Xd_0__inst_mult_8_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_516 ),
	.cout(Xd_0__inst_mult_8_517 ),
	.shareout(Xd_0__inst_mult_8_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_155 (
// Equation(s):
// Xd_0__inst_mult_8_520  = SUM(( (din_a[100] & din_b[105]) ) + ( Xd_0__inst_mult_8_510  ) + ( Xd_0__inst_mult_8_509  ))
// Xd_0__inst_mult_8_521  = CARRY(( (din_a[100] & din_b[105]) ) + ( Xd_0__inst_mult_8_510  ) + ( Xd_0__inst_mult_8_509  ))
// Xd_0__inst_mult_8_522  = SHARE((din_a[100] & din_b[106]))

	.dataa(!din_a[100]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_509 ),
	.sharein(Xd_0__inst_mult_8_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_520 ),
	.cout(Xd_0__inst_mult_8_521 ),
	.shareout(Xd_0__inst_mult_8_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_156 (
// Equation(s):
// Xd_0__inst_mult_8_524  = SUM(( (!din_a[102] & (((din_a[101] & din_b[104])))) # (din_a[102] & (!din_b[103] $ (((!din_a[101]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_514  ) + ( Xd_0__inst_mult_8_513  ))
// Xd_0__inst_mult_8_525  = CARRY(( (!din_a[102] & (((din_a[101] & din_b[104])))) # (din_a[102] & (!din_b[103] $ (((!din_a[101]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_514  ) + ( Xd_0__inst_mult_8_513  ))
// Xd_0__inst_mult_8_526  = SHARE((din_a[102] & (din_b[103] & (din_a[101] & din_b[104]))))

	.dataa(!din_a[102]),
	.datab(!din_b[103]),
	.datac(!din_a[101]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_513 ),
	.sharein(Xd_0__inst_mult_8_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_524 ),
	.cout(Xd_0__inst_mult_8_525 ),
	.shareout(Xd_0__inst_mult_8_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_150 (
// Equation(s):
// Xd_0__inst_mult_9_512  = SUM(( (din_a[116] & din_b[113]) ) + ( Xd_0__inst_mult_9_502  ) + ( Xd_0__inst_mult_9_501  ))
// Xd_0__inst_mult_9_513  = CARRY(( (din_a[116] & din_b[113]) ) + ( Xd_0__inst_mult_9_502  ) + ( Xd_0__inst_mult_9_501  ))
// Xd_0__inst_mult_9_514  = SHARE((din_a[116] & din_b[114]))

	.dataa(!din_a[116]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_501 ),
	.sharein(Xd_0__inst_mult_9_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_512 ),
	.cout(Xd_0__inst_mult_9_513 ),
	.shareout(Xd_0__inst_mult_9_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_151 (
// Equation(s):
// Xd_0__inst_mult_9_516  = SUM(( (din_a[112] & din_b[117]) ) + ( Xd_0__inst_mult_9_506  ) + ( Xd_0__inst_mult_9_505  ))
// Xd_0__inst_mult_9_517  = CARRY(( (din_a[112] & din_b[117]) ) + ( Xd_0__inst_mult_9_506  ) + ( Xd_0__inst_mult_9_505  ))
// Xd_0__inst_mult_9_518  = SHARE((din_a[112] & din_b[118]))

	.dataa(!din_a[112]),
	.datab(!din_b[117]),
	.datac(!din_b[118]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_505 ),
	.sharein(Xd_0__inst_mult_9_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_516 ),
	.cout(Xd_0__inst_mult_9_517 ),
	.shareout(Xd_0__inst_mult_9_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_152 (
// Equation(s):
// Xd_0__inst_mult_9_520  = SUM(( (!din_a[114] & (((din_a[113] & din_b[116])))) # (din_a[114] & (!din_b[115] $ (((!din_a[113]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_510  ) + ( Xd_0__inst_mult_9_509  ))
// Xd_0__inst_mult_9_521  = CARRY(( (!din_a[114] & (((din_a[113] & din_b[116])))) # (din_a[114] & (!din_b[115] $ (((!din_a[113]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_510  ) + ( Xd_0__inst_mult_9_509  ))
// Xd_0__inst_mult_9_522  = SHARE((din_a[114] & (din_b[115] & (din_a[113] & din_b[116]))))

	.dataa(!din_a[114]),
	.datab(!din_b[115]),
	.datac(!din_a[113]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_509 ),
	.sharein(Xd_0__inst_mult_9_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_520 ),
	.cout(Xd_0__inst_mult_9_521 ),
	.shareout(Xd_0__inst_mult_9_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_150 (
// Equation(s):
// Xd_0__inst_mult_6_512  = SUM(( (din_a[80] & din_b[77]) ) + ( Xd_0__inst_mult_6_502  ) + ( Xd_0__inst_mult_6_501  ))
// Xd_0__inst_mult_6_513  = CARRY(( (din_a[80] & din_b[77]) ) + ( Xd_0__inst_mult_6_502  ) + ( Xd_0__inst_mult_6_501  ))
// Xd_0__inst_mult_6_514  = SHARE((din_a[80] & din_b[78]))

	.dataa(!din_a[80]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_501 ),
	.sharein(Xd_0__inst_mult_6_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_512 ),
	.cout(Xd_0__inst_mult_6_513 ),
	.shareout(Xd_0__inst_mult_6_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_151 (
// Equation(s):
// Xd_0__inst_mult_6_516  = SUM(( (din_a[76] & din_b[81]) ) + ( Xd_0__inst_mult_6_506  ) + ( Xd_0__inst_mult_6_505  ))
// Xd_0__inst_mult_6_517  = CARRY(( (din_a[76] & din_b[81]) ) + ( Xd_0__inst_mult_6_506  ) + ( Xd_0__inst_mult_6_505  ))
// Xd_0__inst_mult_6_518  = SHARE((din_a[76] & din_b[82]))

	.dataa(!din_a[76]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_505 ),
	.sharein(Xd_0__inst_mult_6_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_516 ),
	.cout(Xd_0__inst_mult_6_517 ),
	.shareout(Xd_0__inst_mult_6_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_152 (
// Equation(s):
// Xd_0__inst_mult_6_520  = SUM(( (!din_a[78] & (((din_a[77] & din_b[80])))) # (din_a[78] & (!din_b[79] $ (((!din_a[77]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_510  ) + ( Xd_0__inst_mult_6_509  ))
// Xd_0__inst_mult_6_521  = CARRY(( (!din_a[78] & (((din_a[77] & din_b[80])))) # (din_a[78] & (!din_b[79] $ (((!din_a[77]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_510  ) + ( Xd_0__inst_mult_6_509  ))
// Xd_0__inst_mult_6_522  = SHARE((din_a[78] & (din_b[79] & (din_a[77] & din_b[80]))))

	.dataa(!din_a[78]),
	.datab(!din_b[79]),
	.datac(!din_a[77]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_509 ),
	.sharein(Xd_0__inst_mult_6_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_520 ),
	.cout(Xd_0__inst_mult_6_521 ),
	.shareout(Xd_0__inst_mult_6_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_148 (
// Equation(s):
// Xd_0__inst_mult_7_504  = SUM(( (din_a[93] & din_b[88]) ) + ( Xd_0__inst_mult_7_490  ) + ( Xd_0__inst_mult_7_489  ))
// Xd_0__inst_mult_7_505  = CARRY(( (din_a[93] & din_b[88]) ) + ( Xd_0__inst_mult_7_490  ) + ( Xd_0__inst_mult_7_489  ))
// Xd_0__inst_mult_7_506  = SHARE(GND)

	.dataa(!din_a[93]),
	.datab(!din_b[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_489 ),
	.sharein(Xd_0__inst_mult_7_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_504 ),
	.cout(Xd_0__inst_mult_7_505 ),
	.shareout(Xd_0__inst_mult_7_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_149 (
// Equation(s):
// Xd_0__inst_mult_7_508  = SUM(( (din_a[92] & din_b[89]) ) + ( Xd_0__inst_mult_7_494  ) + ( Xd_0__inst_mult_7_493  ))
// Xd_0__inst_mult_7_509  = CARRY(( (din_a[92] & din_b[89]) ) + ( Xd_0__inst_mult_7_494  ) + ( Xd_0__inst_mult_7_493  ))
// Xd_0__inst_mult_7_510  = SHARE((din_a[92] & din_b[90]))

	.dataa(!din_a[92]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_493 ),
	.sharein(Xd_0__inst_mult_7_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_508 ),
	.cout(Xd_0__inst_mult_7_509 ),
	.shareout(Xd_0__inst_mult_7_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_150 (
// Equation(s):
// Xd_0__inst_mult_7_512  = SUM(( (din_a[88] & din_b[93]) ) + ( Xd_0__inst_mult_7_498  ) + ( Xd_0__inst_mult_7_497  ))
// Xd_0__inst_mult_7_513  = CARRY(( (din_a[88] & din_b[93]) ) + ( Xd_0__inst_mult_7_498  ) + ( Xd_0__inst_mult_7_497  ))
// Xd_0__inst_mult_7_514  = SHARE((din_a[88] & din_b[94]))

	.dataa(!din_a[88]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_497 ),
	.sharein(Xd_0__inst_mult_7_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_512 ),
	.cout(Xd_0__inst_mult_7_513 ),
	.shareout(Xd_0__inst_mult_7_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_151 (
// Equation(s):
// Xd_0__inst_mult_7_516  = SUM(( (!din_a[90] & (((din_a[89] & din_b[92])))) # (din_a[90] & (!din_b[91] $ (((!din_a[89]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_502  ) + ( Xd_0__inst_mult_7_501  ))
// Xd_0__inst_mult_7_517  = CARRY(( (!din_a[90] & (((din_a[89] & din_b[92])))) # (din_a[90] & (!din_b[91] $ (((!din_a[89]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_502  ) + ( Xd_0__inst_mult_7_501  ))
// Xd_0__inst_mult_7_518  = SHARE((din_a[90] & (din_b[91] & (din_a[89] & din_b[92]))))

	.dataa(!din_a[90]),
	.datab(!din_b[91]),
	.datac(!din_a[89]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_501 ),
	.sharein(Xd_0__inst_mult_7_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_516 ),
	.cout(Xd_0__inst_mult_7_517 ),
	.shareout(Xd_0__inst_mult_7_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_159 (
// Equation(s):
// Xd_0__inst_mult_4_536  = SUM(( (din_a[57] & din_b[52]) ) + ( Xd_0__inst_mult_4_526  ) + ( Xd_0__inst_mult_4_525  ))
// Xd_0__inst_mult_4_537  = CARRY(( (din_a[57] & din_b[52]) ) + ( Xd_0__inst_mult_4_526  ) + ( Xd_0__inst_mult_4_525  ))
// Xd_0__inst_mult_4_538  = SHARE(GND)

	.dataa(!din_a[57]),
	.datab(!din_b[52]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_525 ),
	.sharein(Xd_0__inst_mult_4_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_536 ),
	.cout(Xd_0__inst_mult_4_537 ),
	.shareout(Xd_0__inst_mult_4_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_160 (
// Equation(s):
// Xd_0__inst_mult_4_540  = SUM(( (din_a[56] & din_b[53]) ) + ( Xd_0__inst_mult_4_530  ) + ( Xd_0__inst_mult_4_529  ))
// Xd_0__inst_mult_4_541  = CARRY(( (din_a[56] & din_b[53]) ) + ( Xd_0__inst_mult_4_530  ) + ( Xd_0__inst_mult_4_529  ))
// Xd_0__inst_mult_4_542  = SHARE((din_a[56] & din_b[54]))

	.dataa(!din_a[56]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_529 ),
	.sharein(Xd_0__inst_mult_4_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_540 ),
	.cout(Xd_0__inst_mult_4_541 ),
	.shareout(Xd_0__inst_mult_4_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_161 (
// Equation(s):
// Xd_0__inst_mult_4_544  = SUM(( (!din_a[54] & (((din_a[53] & din_b[56])))) # (din_a[54] & (!din_b[55] $ (((!din_a[53]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_534  ) + ( Xd_0__inst_mult_4_533  ))
// Xd_0__inst_mult_4_545  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[56])))) # (din_a[54] & (!din_b[55] $ (((!din_a[53]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_534  ) + ( Xd_0__inst_mult_4_533  ))
// Xd_0__inst_mult_4_546  = SHARE((din_a[54] & (din_b[55] & (din_a[53] & din_b[56]))))

	.dataa(!din_a[54]),
	.datab(!din_b[55]),
	.datac(!din_a[53]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_533 ),
	.sharein(Xd_0__inst_mult_4_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_544 ),
	.cout(Xd_0__inst_mult_4_545 ),
	.shareout(Xd_0__inst_mult_4_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_148 (
// Equation(s):
// Xd_0__inst_mult_5_504  = SUM(( (din_a[69] & din_b[64]) ) + ( Xd_0__inst_mult_5_490  ) + ( Xd_0__inst_mult_5_489  ))
// Xd_0__inst_mult_5_505  = CARRY(( (din_a[69] & din_b[64]) ) + ( Xd_0__inst_mult_5_490  ) + ( Xd_0__inst_mult_5_489  ))
// Xd_0__inst_mult_5_506  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[64]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_489 ),
	.sharein(Xd_0__inst_mult_5_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_504 ),
	.cout(Xd_0__inst_mult_5_505 ),
	.shareout(Xd_0__inst_mult_5_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_149 (
// Equation(s):
// Xd_0__inst_mult_5_508  = SUM(( (din_a[68] & din_b[65]) ) + ( Xd_0__inst_mult_5_494  ) + ( Xd_0__inst_mult_5_493  ))
// Xd_0__inst_mult_5_509  = CARRY(( (din_a[68] & din_b[65]) ) + ( Xd_0__inst_mult_5_494  ) + ( Xd_0__inst_mult_5_493  ))
// Xd_0__inst_mult_5_510  = SHARE((din_a[68] & din_b[66]))

	.dataa(!din_a[68]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_493 ),
	.sharein(Xd_0__inst_mult_5_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_508 ),
	.cout(Xd_0__inst_mult_5_509 ),
	.shareout(Xd_0__inst_mult_5_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_150 (
// Equation(s):
// Xd_0__inst_mult_5_512  = SUM(( (din_a[64] & din_b[69]) ) + ( Xd_0__inst_mult_5_498  ) + ( Xd_0__inst_mult_5_497  ))
// Xd_0__inst_mult_5_513  = CARRY(( (din_a[64] & din_b[69]) ) + ( Xd_0__inst_mult_5_498  ) + ( Xd_0__inst_mult_5_497  ))
// Xd_0__inst_mult_5_514  = SHARE((din_a[64] & din_b[70]))

	.dataa(!din_a[64]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_497 ),
	.sharein(Xd_0__inst_mult_5_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_512 ),
	.cout(Xd_0__inst_mult_5_513 ),
	.shareout(Xd_0__inst_mult_5_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_151 (
// Equation(s):
// Xd_0__inst_mult_5_516  = SUM(( (!din_a[66] & (((din_a[65] & din_b[68])))) # (din_a[66] & (!din_b[67] $ (((!din_a[65]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_502  ) + ( Xd_0__inst_mult_5_501  ))
// Xd_0__inst_mult_5_517  = CARRY(( (!din_a[66] & (((din_a[65] & din_b[68])))) # (din_a[66] & (!din_b[67] $ (((!din_a[65]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_502  ) + ( Xd_0__inst_mult_5_501  ))
// Xd_0__inst_mult_5_518  = SHARE((din_a[66] & (din_b[67] & (din_a[65] & din_b[68]))))

	.dataa(!din_a[66]),
	.datab(!din_b[67]),
	.datac(!din_a[65]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_501 ),
	.sharein(Xd_0__inst_mult_5_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_516 ),
	.cout(Xd_0__inst_mult_5_517 ),
	.shareout(Xd_0__inst_mult_5_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_152 (
// Equation(s):
// Xd_0__inst_mult_2_508  = SUM(( (din_a[33] & din_b[28]) ) + ( Xd_0__inst_mult_2_494  ) + ( Xd_0__inst_mult_2_493  ))
// Xd_0__inst_mult_2_509  = CARRY(( (din_a[33] & din_b[28]) ) + ( Xd_0__inst_mult_2_494  ) + ( Xd_0__inst_mult_2_493  ))
// Xd_0__inst_mult_2_510  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_493 ),
	.sharein(Xd_0__inst_mult_2_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_508 ),
	.cout(Xd_0__inst_mult_2_509 ),
	.shareout(Xd_0__inst_mult_2_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_153 (
// Equation(s):
// Xd_0__inst_mult_2_512  = SUM(( (din_a[32] & din_b[29]) ) + ( Xd_0__inst_mult_2_498  ) + ( Xd_0__inst_mult_2_497  ))
// Xd_0__inst_mult_2_513  = CARRY(( (din_a[32] & din_b[29]) ) + ( Xd_0__inst_mult_2_498  ) + ( Xd_0__inst_mult_2_497  ))
// Xd_0__inst_mult_2_514  = SHARE((din_a[32] & din_b[30]))

	.dataa(!din_a[32]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_497 ),
	.sharein(Xd_0__inst_mult_2_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_512 ),
	.cout(Xd_0__inst_mult_2_513 ),
	.shareout(Xd_0__inst_mult_2_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_154 (
// Equation(s):
// Xd_0__inst_mult_2_516  = SUM(( (din_a[28] & din_b[33]) ) + ( Xd_0__inst_mult_2_502  ) + ( Xd_0__inst_mult_2_501  ))
// Xd_0__inst_mult_2_517  = CARRY(( (din_a[28] & din_b[33]) ) + ( Xd_0__inst_mult_2_502  ) + ( Xd_0__inst_mult_2_501  ))
// Xd_0__inst_mult_2_518  = SHARE((din_a[28] & din_b[34]))

	.dataa(!din_a[28]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_501 ),
	.sharein(Xd_0__inst_mult_2_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_516 ),
	.cout(Xd_0__inst_mult_2_517 ),
	.shareout(Xd_0__inst_mult_2_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_155 (
// Equation(s):
// Xd_0__inst_mult_2_520  = SUM(( (!din_a[30] & (((din_a[29] & din_b[32])))) # (din_a[30] & (!din_b[31] $ (((!din_a[29]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_506  ) + ( Xd_0__inst_mult_2_505  ))
// Xd_0__inst_mult_2_521  = CARRY(( (!din_a[30] & (((din_a[29] & din_b[32])))) # (din_a[30] & (!din_b[31] $ (((!din_a[29]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_506  ) + ( Xd_0__inst_mult_2_505  ))
// Xd_0__inst_mult_2_522  = SHARE((din_a[30] & (din_b[31] & (din_a[29] & din_b[32]))))

	.dataa(!din_a[30]),
	.datab(!din_b[31]),
	.datac(!din_a[29]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_505 ),
	.sharein(Xd_0__inst_mult_2_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_520 ),
	.cout(Xd_0__inst_mult_2_521 ),
	.shareout(Xd_0__inst_mult_2_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_148 (
// Equation(s):
// Xd_0__inst_mult_3_504  = SUM(( (din_a[45] & din_b[40]) ) + ( Xd_0__inst_mult_3_490  ) + ( Xd_0__inst_mult_3_489  ))
// Xd_0__inst_mult_3_505  = CARRY(( (din_a[45] & din_b[40]) ) + ( Xd_0__inst_mult_3_490  ) + ( Xd_0__inst_mult_3_489  ))
// Xd_0__inst_mult_3_506  = SHARE(GND)

	.dataa(!din_a[45]),
	.datab(!din_b[40]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_489 ),
	.sharein(Xd_0__inst_mult_3_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_504 ),
	.cout(Xd_0__inst_mult_3_505 ),
	.shareout(Xd_0__inst_mult_3_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_149 (
// Equation(s):
// Xd_0__inst_mult_3_508  = SUM(( (din_a[44] & din_b[41]) ) + ( Xd_0__inst_mult_3_494  ) + ( Xd_0__inst_mult_3_493  ))
// Xd_0__inst_mult_3_509  = CARRY(( (din_a[44] & din_b[41]) ) + ( Xd_0__inst_mult_3_494  ) + ( Xd_0__inst_mult_3_493  ))
// Xd_0__inst_mult_3_510  = SHARE((din_a[44] & din_b[42]))

	.dataa(!din_a[44]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_493 ),
	.sharein(Xd_0__inst_mult_3_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_508 ),
	.cout(Xd_0__inst_mult_3_509 ),
	.shareout(Xd_0__inst_mult_3_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_150 (
// Equation(s):
// Xd_0__inst_mult_3_512  = SUM(( (din_a[40] & din_b[45]) ) + ( Xd_0__inst_mult_3_498  ) + ( Xd_0__inst_mult_3_497  ))
// Xd_0__inst_mult_3_513  = CARRY(( (din_a[40] & din_b[45]) ) + ( Xd_0__inst_mult_3_498  ) + ( Xd_0__inst_mult_3_497  ))
// Xd_0__inst_mult_3_514  = SHARE((din_a[40] & din_b[46]))

	.dataa(!din_a[40]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_497 ),
	.sharein(Xd_0__inst_mult_3_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_512 ),
	.cout(Xd_0__inst_mult_3_513 ),
	.shareout(Xd_0__inst_mult_3_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_151 (
// Equation(s):
// Xd_0__inst_mult_3_516  = SUM(( (!din_a[42] & (((din_a[41] & din_b[44])))) # (din_a[42] & (!din_b[43] $ (((!din_a[41]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_502  ) + ( Xd_0__inst_mult_3_501  ))
// Xd_0__inst_mult_3_517  = CARRY(( (!din_a[42] & (((din_a[41] & din_b[44])))) # (din_a[42] & (!din_b[43] $ (((!din_a[41]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_502  ) + ( Xd_0__inst_mult_3_501  ))
// Xd_0__inst_mult_3_518  = SHARE((din_a[42] & (din_b[43] & (din_a[41] & din_b[44]))))

	.dataa(!din_a[42]),
	.datab(!din_b[43]),
	.datac(!din_a[41]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_501 ),
	.sharein(Xd_0__inst_mult_3_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_516 ),
	.cout(Xd_0__inst_mult_3_517 ),
	.shareout(Xd_0__inst_mult_3_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_152 (
// Equation(s):
// Xd_0__inst_mult_0_508  = SUM(( (din_a[9] & din_b[4]) ) + ( Xd_0__inst_mult_0_494  ) + ( Xd_0__inst_mult_0_493  ))
// Xd_0__inst_mult_0_509  = CARRY(( (din_a[9] & din_b[4]) ) + ( Xd_0__inst_mult_0_494  ) + ( Xd_0__inst_mult_0_493  ))
// Xd_0__inst_mult_0_510  = SHARE(GND)

	.dataa(!din_a[9]),
	.datab(!din_b[4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_493 ),
	.sharein(Xd_0__inst_mult_0_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_508 ),
	.cout(Xd_0__inst_mult_0_509 ),
	.shareout(Xd_0__inst_mult_0_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_153 (
// Equation(s):
// Xd_0__inst_mult_0_512  = SUM(( (din_a[8] & din_b[5]) ) + ( Xd_0__inst_mult_0_498  ) + ( Xd_0__inst_mult_0_497  ))
// Xd_0__inst_mult_0_513  = CARRY(( (din_a[8] & din_b[5]) ) + ( Xd_0__inst_mult_0_498  ) + ( Xd_0__inst_mult_0_497  ))
// Xd_0__inst_mult_0_514  = SHARE((din_a[8] & din_b[6]))

	.dataa(!din_a[8]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_497 ),
	.sharein(Xd_0__inst_mult_0_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_512 ),
	.cout(Xd_0__inst_mult_0_513 ),
	.shareout(Xd_0__inst_mult_0_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_154 (
// Equation(s):
// Xd_0__inst_mult_0_516  = SUM(( (din_a[4] & din_b[9]) ) + ( Xd_0__inst_mult_0_502  ) + ( Xd_0__inst_mult_0_501  ))
// Xd_0__inst_mult_0_517  = CARRY(( (din_a[4] & din_b[9]) ) + ( Xd_0__inst_mult_0_502  ) + ( Xd_0__inst_mult_0_501  ))
// Xd_0__inst_mult_0_518  = SHARE((din_a[4] & din_b[10]))

	.dataa(!din_a[4]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_501 ),
	.sharein(Xd_0__inst_mult_0_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_516 ),
	.cout(Xd_0__inst_mult_0_517 ),
	.shareout(Xd_0__inst_mult_0_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_155 (
// Equation(s):
// Xd_0__inst_mult_0_520  = SUM(( (!din_a[6] & (((din_a[5] & din_b[8])))) # (din_a[6] & (!din_b[7] $ (((!din_a[5]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_506  ) + ( Xd_0__inst_mult_0_505  ))
// Xd_0__inst_mult_0_521  = CARRY(( (!din_a[6] & (((din_a[5] & din_b[8])))) # (din_a[6] & (!din_b[7] $ (((!din_a[5]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_506  ) + ( Xd_0__inst_mult_0_505  ))
// Xd_0__inst_mult_0_522  = SHARE((din_a[6] & (din_b[7] & (din_a[5] & din_b[8]))))

	.dataa(!din_a[6]),
	.datab(!din_b[7]),
	.datac(!din_a[5]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_505 ),
	.sharein(Xd_0__inst_mult_0_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_520 ),
	.cout(Xd_0__inst_mult_0_521 ),
	.shareout(Xd_0__inst_mult_0_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_152 (
// Equation(s):
// Xd_0__inst_mult_1_508  = SUM(( (din_a[21] & din_b[16]) ) + ( Xd_0__inst_mult_1_494  ) + ( Xd_0__inst_mult_1_493  ))
// Xd_0__inst_mult_1_509  = CARRY(( (din_a[21] & din_b[16]) ) + ( Xd_0__inst_mult_1_494  ) + ( Xd_0__inst_mult_1_493  ))
// Xd_0__inst_mult_1_510  = SHARE(GND)

	.dataa(!din_a[21]),
	.datab(!din_b[16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_493 ),
	.sharein(Xd_0__inst_mult_1_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_508 ),
	.cout(Xd_0__inst_mult_1_509 ),
	.shareout(Xd_0__inst_mult_1_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_153 (
// Equation(s):
// Xd_0__inst_mult_1_512  = SUM(( (din_a[20] & din_b[17]) ) + ( Xd_0__inst_mult_1_498  ) + ( Xd_0__inst_mult_1_497  ))
// Xd_0__inst_mult_1_513  = CARRY(( (din_a[20] & din_b[17]) ) + ( Xd_0__inst_mult_1_498  ) + ( Xd_0__inst_mult_1_497  ))
// Xd_0__inst_mult_1_514  = SHARE((din_a[20] & din_b[18]))

	.dataa(!din_a[20]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_497 ),
	.sharein(Xd_0__inst_mult_1_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_512 ),
	.cout(Xd_0__inst_mult_1_513 ),
	.shareout(Xd_0__inst_mult_1_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_154 (
// Equation(s):
// Xd_0__inst_mult_1_516  = SUM(( (din_a[16] & din_b[21]) ) + ( Xd_0__inst_mult_1_502  ) + ( Xd_0__inst_mult_1_501  ))
// Xd_0__inst_mult_1_517  = CARRY(( (din_a[16] & din_b[21]) ) + ( Xd_0__inst_mult_1_502  ) + ( Xd_0__inst_mult_1_501  ))
// Xd_0__inst_mult_1_518  = SHARE((din_a[16] & din_b[22]))

	.dataa(!din_a[16]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_501 ),
	.sharein(Xd_0__inst_mult_1_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_516 ),
	.cout(Xd_0__inst_mult_1_517 ),
	.shareout(Xd_0__inst_mult_1_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_155 (
// Equation(s):
// Xd_0__inst_mult_1_520  = SUM(( (!din_a[18] & (((din_a[17] & din_b[20])))) # (din_a[18] & (!din_b[19] $ (((!din_a[17]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_506  ) + ( Xd_0__inst_mult_1_505  ))
// Xd_0__inst_mult_1_521  = CARRY(( (!din_a[18] & (((din_a[17] & din_b[20])))) # (din_a[18] & (!din_b[19] $ (((!din_a[17]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_506  ) + ( Xd_0__inst_mult_1_505  ))
// Xd_0__inst_mult_1_522  = SHARE((din_a[18] & (din_b[19] & (din_a[17] & din_b[20]))))

	.dataa(!din_a[18]),
	.datab(!din_b[19]),
	.datac(!din_a[17]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_505 ),
	.sharein(Xd_0__inst_mult_1_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_520 ),
	.cout(Xd_0__inst_mult_1_521 ),
	.shareout(Xd_0__inst_mult_1_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_159 (
// Equation(s):
// Xd_0__inst_mult_12_548  = SUM(( (din_a[153] & din_b[149]) ) + ( Xd_0__inst_mult_12_542  ) + ( Xd_0__inst_mult_12_541  ))
// Xd_0__inst_mult_12_549  = CARRY(( (din_a[153] & din_b[149]) ) + ( Xd_0__inst_mult_12_542  ) + ( Xd_0__inst_mult_12_541  ))
// Xd_0__inst_mult_12_550  = SHARE((din_a[153] & din_b[150]))

	.dataa(!din_a[153]),
	.datab(!din_b[149]),
	.datac(!din_b[150]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_541 ),
	.sharein(Xd_0__inst_mult_12_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_548 ),
	.cout(Xd_0__inst_mult_12_549 ),
	.shareout(Xd_0__inst_mult_12_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_160 (
// Equation(s):
// Xd_0__inst_mult_12_552  = SUM(( (!din_a[151] & (((din_a[150] & din_b[152])))) # (din_a[151] & (!din_b[151] $ (((!din_a[150]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_546  ) + ( Xd_0__inst_mult_12_545  ))
// Xd_0__inst_mult_12_553  = CARRY(( (!din_a[151] & (((din_a[150] & din_b[152])))) # (din_a[151] & (!din_b[151] $ (((!din_a[150]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_12_546  ) + ( Xd_0__inst_mult_12_545  ))
// Xd_0__inst_mult_12_554  = SHARE((din_a[151] & (din_b[151] & (din_a[150] & din_b[152]))))

	.dataa(!din_a[151]),
	.datab(!din_b[151]),
	.datac(!din_a[150]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_545 ),
	.sharein(Xd_0__inst_mult_12_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_552 ),
	.cout(Xd_0__inst_mult_12_553 ),
	.shareout(Xd_0__inst_mult_12_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_157 (
// Equation(s):
// Xd_0__inst_mult_13_528  = SUM(( (din_a[165] & din_b[161]) ) + ( Xd_0__inst_mult_13_518  ) + ( Xd_0__inst_mult_13_517  ))
// Xd_0__inst_mult_13_529  = CARRY(( (din_a[165] & din_b[161]) ) + ( Xd_0__inst_mult_13_518  ) + ( Xd_0__inst_mult_13_517  ))
// Xd_0__inst_mult_13_530  = SHARE((din_a[165] & din_b[162]))

	.dataa(!din_a[165]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_517 ),
	.sharein(Xd_0__inst_mult_13_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_528 ),
	.cout(Xd_0__inst_mult_13_529 ),
	.shareout(Xd_0__inst_mult_13_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_158 (
// Equation(s):
// Xd_0__inst_mult_13_532  = SUM(( (din_a[161] & din_b[165]) ) + ( Xd_0__inst_mult_13_522  ) + ( Xd_0__inst_mult_13_521  ))
// Xd_0__inst_mult_13_533  = CARRY(( (din_a[161] & din_b[165]) ) + ( Xd_0__inst_mult_13_522  ) + ( Xd_0__inst_mult_13_521  ))
// Xd_0__inst_mult_13_534  = SHARE((din_a[161] & din_b[166]))

	.dataa(!din_a[161]),
	.datab(!din_b[165]),
	.datac(!din_b[166]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_521 ),
	.sharein(Xd_0__inst_mult_13_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_532 ),
	.cout(Xd_0__inst_mult_13_533 ),
	.shareout(Xd_0__inst_mult_13_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_159 (
// Equation(s):
// Xd_0__inst_mult_13_536  = SUM(( (!din_a[163] & (((din_a[162] & din_b[164])))) # (din_a[163] & (!din_b[163] $ (((!din_a[162]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_526  ) + ( Xd_0__inst_mult_13_525  ))
// Xd_0__inst_mult_13_537  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[164])))) # (din_a[163] & (!din_b[163] $ (((!din_a[162]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_13_526  ) + ( Xd_0__inst_mult_13_525  ))
// Xd_0__inst_mult_13_538  = SHARE((din_a[163] & (din_b[163] & (din_a[162] & din_b[164]))))

	.dataa(!din_a[163]),
	.datab(!din_b[163]),
	.datac(!din_a[162]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_525 ),
	.sharein(Xd_0__inst_mult_13_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_536 ),
	.cout(Xd_0__inst_mult_13_537 ),
	.shareout(Xd_0__inst_mult_13_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_157 (
// Equation(s):
// Xd_0__inst_mult_14_528  = SUM(( (din_a[177] & din_b[173]) ) + ( Xd_0__inst_mult_14_518  ) + ( Xd_0__inst_mult_14_517  ))
// Xd_0__inst_mult_14_529  = CARRY(( (din_a[177] & din_b[173]) ) + ( Xd_0__inst_mult_14_518  ) + ( Xd_0__inst_mult_14_517  ))
// Xd_0__inst_mult_14_530  = SHARE((din_a[177] & din_b[174]))

	.dataa(!din_a[177]),
	.datab(!din_b[173]),
	.datac(!din_b[174]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_517 ),
	.sharein(Xd_0__inst_mult_14_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_528 ),
	.cout(Xd_0__inst_mult_14_529 ),
	.shareout(Xd_0__inst_mult_14_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_158 (
// Equation(s):
// Xd_0__inst_mult_14_532  = SUM(( (din_a[173] & din_b[177]) ) + ( Xd_0__inst_mult_14_522  ) + ( Xd_0__inst_mult_14_521  ))
// Xd_0__inst_mult_14_533  = CARRY(( (din_a[173] & din_b[177]) ) + ( Xd_0__inst_mult_14_522  ) + ( Xd_0__inst_mult_14_521  ))
// Xd_0__inst_mult_14_534  = SHARE((din_a[173] & din_b[178]))

	.dataa(!din_a[173]),
	.datab(!din_b[177]),
	.datac(!din_b[178]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_521 ),
	.sharein(Xd_0__inst_mult_14_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_532 ),
	.cout(Xd_0__inst_mult_14_533 ),
	.shareout(Xd_0__inst_mult_14_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_159 (
// Equation(s):
// Xd_0__inst_mult_14_536  = SUM(( (!din_a[175] & (((din_a[174] & din_b[176])))) # (din_a[175] & (!din_b[175] $ (((!din_a[174]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_526  ) + ( Xd_0__inst_mult_14_525  ))
// Xd_0__inst_mult_14_537  = CARRY(( (!din_a[175] & (((din_a[174] & din_b[176])))) # (din_a[175] & (!din_b[175] $ (((!din_a[174]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_14_526  ) + ( Xd_0__inst_mult_14_525  ))
// Xd_0__inst_mult_14_538  = SHARE((din_a[175] & (din_b[175] & (din_a[174] & din_b[176]))))

	.dataa(!din_a[175]),
	.datab(!din_b[175]),
	.datac(!din_a[174]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_525 ),
	.sharein(Xd_0__inst_mult_14_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_536 ),
	.cout(Xd_0__inst_mult_14_537 ),
	.shareout(Xd_0__inst_mult_14_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_163 (
// Equation(s):
// Xd_0__inst_mult_15_552  = SUM(( (din_a[189] & din_b[185]) ) + ( Xd_0__inst_mult_15_546  ) + ( Xd_0__inst_mult_15_545  ))
// Xd_0__inst_mult_15_553  = CARRY(( (din_a[189] & din_b[185]) ) + ( Xd_0__inst_mult_15_546  ) + ( Xd_0__inst_mult_15_545  ))
// Xd_0__inst_mult_15_554  = SHARE((din_a[189] & din_b[186]))

	.dataa(!din_a[189]),
	.datab(!din_b[185]),
	.datac(!din_b[186]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_545 ),
	.sharein(Xd_0__inst_mult_15_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_552 ),
	.cout(Xd_0__inst_mult_15_553 ),
	.shareout(Xd_0__inst_mult_15_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_164 (
// Equation(s):
// Xd_0__inst_mult_15_556  = SUM(( (!din_a[187] & (((din_a[186] & din_b[188])))) # (din_a[187] & (!din_b[187] $ (((!din_a[186]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_550  ) + ( Xd_0__inst_mult_15_549  ))
// Xd_0__inst_mult_15_557  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[188])))) # (din_a[187] & (!din_b[187] $ (((!din_a[186]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_15_550  ) + ( Xd_0__inst_mult_15_549  ))
// Xd_0__inst_mult_15_558  = SHARE((din_a[187] & (din_b[187] & (din_a[186] & din_b[188]))))

	.dataa(!din_a[187]),
	.datab(!din_b[187]),
	.datac(!din_a[186]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_549 ),
	.sharein(Xd_0__inst_mult_15_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_556 ),
	.cout(Xd_0__inst_mult_15_557 ),
	.shareout(Xd_0__inst_mult_15_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_153 (
// Equation(s):
// Xd_0__inst_mult_10_524  = SUM(( (din_a[129] & din_b[125]) ) + ( Xd_0__inst_mult_10_514  ) + ( Xd_0__inst_mult_10_513  ))
// Xd_0__inst_mult_10_525  = CARRY(( (din_a[129] & din_b[125]) ) + ( Xd_0__inst_mult_10_514  ) + ( Xd_0__inst_mult_10_513  ))
// Xd_0__inst_mult_10_526  = SHARE((din_a[129] & din_b[126]))

	.dataa(!din_a[129]),
	.datab(!din_b[125]),
	.datac(!din_b[126]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_513 ),
	.sharein(Xd_0__inst_mult_10_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_524 ),
	.cout(Xd_0__inst_mult_10_525 ),
	.shareout(Xd_0__inst_mult_10_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_154 (
// Equation(s):
// Xd_0__inst_mult_10_528  = SUM(( (din_a[125] & din_b[129]) ) + ( Xd_0__inst_mult_10_518  ) + ( Xd_0__inst_mult_10_517  ))
// Xd_0__inst_mult_10_529  = CARRY(( (din_a[125] & din_b[129]) ) + ( Xd_0__inst_mult_10_518  ) + ( Xd_0__inst_mult_10_517  ))
// Xd_0__inst_mult_10_530  = SHARE((din_a[125] & din_b[130]))

	.dataa(!din_a[125]),
	.datab(!din_b[129]),
	.datac(!din_b[130]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_517 ),
	.sharein(Xd_0__inst_mult_10_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_528 ),
	.cout(Xd_0__inst_mult_10_529 ),
	.shareout(Xd_0__inst_mult_10_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_155 (
// Equation(s):
// Xd_0__inst_mult_10_532  = SUM(( (!din_a[127] & (((din_a[126] & din_b[128])))) # (din_a[127] & (!din_b[127] $ (((!din_a[126]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_522  ) + ( Xd_0__inst_mult_10_521  ))
// Xd_0__inst_mult_10_533  = CARRY(( (!din_a[127] & (((din_a[126] & din_b[128])))) # (din_a[127] & (!din_b[127] $ (((!din_a[126]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_10_522  ) + ( Xd_0__inst_mult_10_521  ))
// Xd_0__inst_mult_10_534  = SHARE((din_a[127] & (din_b[127] & (din_a[126] & din_b[128]))))

	.dataa(!din_a[127]),
	.datab(!din_b[127]),
	.datac(!din_a[126]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_521 ),
	.sharein(Xd_0__inst_mult_10_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_532 ),
	.cout(Xd_0__inst_mult_10_533 ),
	.shareout(Xd_0__inst_mult_10_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_157 (
// Equation(s):
// Xd_0__inst_mult_11_528  = SUM(( (din_a[141] & din_b[137]) ) + ( Xd_0__inst_mult_11_518  ) + ( Xd_0__inst_mult_11_517  ))
// Xd_0__inst_mult_11_529  = CARRY(( (din_a[141] & din_b[137]) ) + ( Xd_0__inst_mult_11_518  ) + ( Xd_0__inst_mult_11_517  ))
// Xd_0__inst_mult_11_530  = SHARE((din_a[141] & din_b[138]))

	.dataa(!din_a[141]),
	.datab(!din_b[137]),
	.datac(!din_b[138]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_517 ),
	.sharein(Xd_0__inst_mult_11_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_528 ),
	.cout(Xd_0__inst_mult_11_529 ),
	.shareout(Xd_0__inst_mult_11_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_158 (
// Equation(s):
// Xd_0__inst_mult_11_532  = SUM(( (din_a[137] & din_b[141]) ) + ( Xd_0__inst_mult_11_522  ) + ( Xd_0__inst_mult_11_521  ))
// Xd_0__inst_mult_11_533  = CARRY(( (din_a[137] & din_b[141]) ) + ( Xd_0__inst_mult_11_522  ) + ( Xd_0__inst_mult_11_521  ))
// Xd_0__inst_mult_11_534  = SHARE((din_a[137] & din_b[142]))

	.dataa(!din_a[137]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_521 ),
	.sharein(Xd_0__inst_mult_11_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_532 ),
	.cout(Xd_0__inst_mult_11_533 ),
	.shareout(Xd_0__inst_mult_11_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_159 (
// Equation(s):
// Xd_0__inst_mult_11_536  = SUM(( (!din_a[139] & (((din_a[138] & din_b[140])))) # (din_a[139] & (!din_b[139] $ (((!din_a[138]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_526  ) + ( Xd_0__inst_mult_11_525  ))
// Xd_0__inst_mult_11_537  = CARRY(( (!din_a[139] & (((din_a[138] & din_b[140])))) # (din_a[139] & (!din_b[139] $ (((!din_a[138]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_11_526  ) + ( Xd_0__inst_mult_11_525  ))
// Xd_0__inst_mult_11_538  = SHARE((din_a[139] & (din_b[139] & (din_a[138] & din_b[140]))))

	.dataa(!din_a[139]),
	.datab(!din_b[139]),
	.datac(!din_a[138]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_525 ),
	.sharein(Xd_0__inst_mult_11_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_536 ),
	.cout(Xd_0__inst_mult_11_537 ),
	.shareout(Xd_0__inst_mult_11_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_157 (
// Equation(s):
// Xd_0__inst_mult_8_528  = SUM(( (din_a[105] & din_b[101]) ) + ( Xd_0__inst_mult_8_518  ) + ( Xd_0__inst_mult_8_517  ))
// Xd_0__inst_mult_8_529  = CARRY(( (din_a[105] & din_b[101]) ) + ( Xd_0__inst_mult_8_518  ) + ( Xd_0__inst_mult_8_517  ))
// Xd_0__inst_mult_8_530  = SHARE((din_a[105] & din_b[102]))

	.dataa(!din_a[105]),
	.datab(!din_b[101]),
	.datac(!din_b[102]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_517 ),
	.sharein(Xd_0__inst_mult_8_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_528 ),
	.cout(Xd_0__inst_mult_8_529 ),
	.shareout(Xd_0__inst_mult_8_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_158 (
// Equation(s):
// Xd_0__inst_mult_8_532  = SUM(( (din_a[101] & din_b[105]) ) + ( Xd_0__inst_mult_8_522  ) + ( Xd_0__inst_mult_8_521  ))
// Xd_0__inst_mult_8_533  = CARRY(( (din_a[101] & din_b[105]) ) + ( Xd_0__inst_mult_8_522  ) + ( Xd_0__inst_mult_8_521  ))
// Xd_0__inst_mult_8_534  = SHARE((din_a[101] & din_b[106]))

	.dataa(!din_a[101]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_521 ),
	.sharein(Xd_0__inst_mult_8_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_532 ),
	.cout(Xd_0__inst_mult_8_533 ),
	.shareout(Xd_0__inst_mult_8_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_159 (
// Equation(s):
// Xd_0__inst_mult_8_536  = SUM(( (!din_a[103] & (((din_a[102] & din_b[104])))) # (din_a[103] & (!din_b[103] $ (((!din_a[102]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_526  ) + ( Xd_0__inst_mult_8_525  ))
// Xd_0__inst_mult_8_537  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[104])))) # (din_a[103] & (!din_b[103] $ (((!din_a[102]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_8_526  ) + ( Xd_0__inst_mult_8_525  ))
// Xd_0__inst_mult_8_538  = SHARE((din_a[103] & (din_b[103] & (din_a[102] & din_b[104]))))

	.dataa(!din_a[103]),
	.datab(!din_b[103]),
	.datac(!din_a[102]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_525 ),
	.sharein(Xd_0__inst_mult_8_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_536 ),
	.cout(Xd_0__inst_mult_8_537 ),
	.shareout(Xd_0__inst_mult_8_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_153 (
// Equation(s):
// Xd_0__inst_mult_9_524  = SUM(( (din_a[117] & din_b[113]) ) + ( Xd_0__inst_mult_9_514  ) + ( Xd_0__inst_mult_9_513  ))
// Xd_0__inst_mult_9_525  = CARRY(( (din_a[117] & din_b[113]) ) + ( Xd_0__inst_mult_9_514  ) + ( Xd_0__inst_mult_9_513  ))
// Xd_0__inst_mult_9_526  = SHARE((din_a[117] & din_b[114]))

	.dataa(!din_a[117]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_513 ),
	.sharein(Xd_0__inst_mult_9_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_524 ),
	.cout(Xd_0__inst_mult_9_525 ),
	.shareout(Xd_0__inst_mult_9_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_154 (
// Equation(s):
// Xd_0__inst_mult_9_528  = SUM(( (din_a[113] & din_b[117]) ) + ( Xd_0__inst_mult_9_518  ) + ( Xd_0__inst_mult_9_517  ))
// Xd_0__inst_mult_9_529  = CARRY(( (din_a[113] & din_b[117]) ) + ( Xd_0__inst_mult_9_518  ) + ( Xd_0__inst_mult_9_517  ))
// Xd_0__inst_mult_9_530  = SHARE((din_a[113] & din_b[118]))

	.dataa(!din_a[113]),
	.datab(!din_b[117]),
	.datac(!din_b[118]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_517 ),
	.sharein(Xd_0__inst_mult_9_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_528 ),
	.cout(Xd_0__inst_mult_9_529 ),
	.shareout(Xd_0__inst_mult_9_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_155 (
// Equation(s):
// Xd_0__inst_mult_9_532  = SUM(( (!din_a[115] & (((din_a[114] & din_b[116])))) # (din_a[115] & (!din_b[115] $ (((!din_a[114]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_522  ) + ( Xd_0__inst_mult_9_521  ))
// Xd_0__inst_mult_9_533  = CARRY(( (!din_a[115] & (((din_a[114] & din_b[116])))) # (din_a[115] & (!din_b[115] $ (((!din_a[114]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_9_522  ) + ( Xd_0__inst_mult_9_521  ))
// Xd_0__inst_mult_9_534  = SHARE((din_a[115] & (din_b[115] & (din_a[114] & din_b[116]))))

	.dataa(!din_a[115]),
	.datab(!din_b[115]),
	.datac(!din_a[114]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_521 ),
	.sharein(Xd_0__inst_mult_9_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_532 ),
	.cout(Xd_0__inst_mult_9_533 ),
	.shareout(Xd_0__inst_mult_9_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_153 (
// Equation(s):
// Xd_0__inst_mult_6_524  = SUM(( (din_a[81] & din_b[77]) ) + ( Xd_0__inst_mult_6_514  ) + ( Xd_0__inst_mult_6_513  ))
// Xd_0__inst_mult_6_525  = CARRY(( (din_a[81] & din_b[77]) ) + ( Xd_0__inst_mult_6_514  ) + ( Xd_0__inst_mult_6_513  ))
// Xd_0__inst_mult_6_526  = SHARE((din_a[81] & din_b[78]))

	.dataa(!din_a[81]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_513 ),
	.sharein(Xd_0__inst_mult_6_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_524 ),
	.cout(Xd_0__inst_mult_6_525 ),
	.shareout(Xd_0__inst_mult_6_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_154 (
// Equation(s):
// Xd_0__inst_mult_6_528  = SUM(( (din_a[77] & din_b[81]) ) + ( Xd_0__inst_mult_6_518  ) + ( Xd_0__inst_mult_6_517  ))
// Xd_0__inst_mult_6_529  = CARRY(( (din_a[77] & din_b[81]) ) + ( Xd_0__inst_mult_6_518  ) + ( Xd_0__inst_mult_6_517  ))
// Xd_0__inst_mult_6_530  = SHARE((din_a[77] & din_b[82]))

	.dataa(!din_a[77]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_517 ),
	.sharein(Xd_0__inst_mult_6_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_528 ),
	.cout(Xd_0__inst_mult_6_529 ),
	.shareout(Xd_0__inst_mult_6_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_155 (
// Equation(s):
// Xd_0__inst_mult_6_532  = SUM(( (!din_a[79] & (((din_a[78] & din_b[80])))) # (din_a[79] & (!din_b[79] $ (((!din_a[78]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_522  ) + ( Xd_0__inst_mult_6_521  ))
// Xd_0__inst_mult_6_533  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[80])))) # (din_a[79] & (!din_b[79] $ (((!din_a[78]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_522  ) + ( Xd_0__inst_mult_6_521  ))
// Xd_0__inst_mult_6_534  = SHARE((din_a[79] & (din_b[79] & (din_a[78] & din_b[80]))))

	.dataa(!din_a[79]),
	.datab(!din_b[79]),
	.datac(!din_a[78]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_521 ),
	.sharein(Xd_0__inst_mult_6_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_532 ),
	.cout(Xd_0__inst_mult_6_533 ),
	.shareout(Xd_0__inst_mult_6_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_152 (
// Equation(s):
// Xd_0__inst_mult_7_520  = SUM(( GND ) + ( Xd_0__inst_mult_7_506  ) + ( Xd_0__inst_mult_7_505  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_505 ),
	.sharein(Xd_0__inst_mult_7_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_520 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_153 (
// Equation(s):
// Xd_0__inst_mult_7_524  = SUM(( (din_a[93] & din_b[89]) ) + ( Xd_0__inst_mult_7_510  ) + ( Xd_0__inst_mult_7_509  ))
// Xd_0__inst_mult_7_525  = CARRY(( (din_a[93] & din_b[89]) ) + ( Xd_0__inst_mult_7_510  ) + ( Xd_0__inst_mult_7_509  ))
// Xd_0__inst_mult_7_526  = SHARE((din_a[93] & din_b[90]))

	.dataa(!din_a[93]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_509 ),
	.sharein(Xd_0__inst_mult_7_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_524 ),
	.cout(Xd_0__inst_mult_7_525 ),
	.shareout(Xd_0__inst_mult_7_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_154 (
// Equation(s):
// Xd_0__inst_mult_7_528  = SUM(( (din_a[89] & din_b[93]) ) + ( Xd_0__inst_mult_7_514  ) + ( Xd_0__inst_mult_7_513  ))
// Xd_0__inst_mult_7_529  = CARRY(( (din_a[89] & din_b[93]) ) + ( Xd_0__inst_mult_7_514  ) + ( Xd_0__inst_mult_7_513  ))
// Xd_0__inst_mult_7_530  = SHARE((din_a[89] & din_b[94]))

	.dataa(!din_a[89]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_513 ),
	.sharein(Xd_0__inst_mult_7_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_528 ),
	.cout(Xd_0__inst_mult_7_529 ),
	.shareout(Xd_0__inst_mult_7_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_155 (
// Equation(s):
// Xd_0__inst_mult_7_532  = SUM(( (!din_a[91] & (((din_a[90] & din_b[92])))) # (din_a[91] & (!din_b[91] $ (((!din_a[90]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_518  ) + ( Xd_0__inst_mult_7_517  ))
// Xd_0__inst_mult_7_533  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[92])))) # (din_a[91] & (!din_b[91] $ (((!din_a[90]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_518  ) + ( Xd_0__inst_mult_7_517  ))
// Xd_0__inst_mult_7_534  = SHARE((din_a[91] & (din_b[91] & (din_a[90] & din_b[92]))))

	.dataa(!din_a[91]),
	.datab(!din_b[91]),
	.datac(!din_a[90]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_517 ),
	.sharein(Xd_0__inst_mult_7_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_532 ),
	.cout(Xd_0__inst_mult_7_533 ),
	.shareout(Xd_0__inst_mult_7_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_162 (
// Equation(s):
// Xd_0__inst_mult_4_548  = SUM(( GND ) + ( Xd_0__inst_mult_4_538  ) + ( Xd_0__inst_mult_4_537  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_537 ),
	.sharein(Xd_0__inst_mult_4_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_548 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_163 (
// Equation(s):
// Xd_0__inst_mult_4_552  = SUM(( (din_a[57] & din_b[53]) ) + ( Xd_0__inst_mult_4_542  ) + ( Xd_0__inst_mult_4_541  ))
// Xd_0__inst_mult_4_553  = CARRY(( (din_a[57] & din_b[53]) ) + ( Xd_0__inst_mult_4_542  ) + ( Xd_0__inst_mult_4_541  ))
// Xd_0__inst_mult_4_554  = SHARE((din_a[57] & din_b[54]))

	.dataa(!din_a[57]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_541 ),
	.sharein(Xd_0__inst_mult_4_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_552 ),
	.cout(Xd_0__inst_mult_4_553 ),
	.shareout(Xd_0__inst_mult_4_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_164 (
// Equation(s):
// Xd_0__inst_mult_4_556  = SUM(( (!din_a[55] & (((din_a[54] & din_b[56])))) # (din_a[55] & (!din_b[55] $ (((!din_a[54]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_546  ) + ( Xd_0__inst_mult_4_545  ))
// Xd_0__inst_mult_4_557  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[56])))) # (din_a[55] & (!din_b[55] $ (((!din_a[54]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_546  ) + ( Xd_0__inst_mult_4_545  ))
// Xd_0__inst_mult_4_558  = SHARE((din_a[55] & (din_b[55] & (din_a[54] & din_b[56]))))

	.dataa(!din_a[55]),
	.datab(!din_b[55]),
	.datac(!din_a[54]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_545 ),
	.sharein(Xd_0__inst_mult_4_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_556 ),
	.cout(Xd_0__inst_mult_4_557 ),
	.shareout(Xd_0__inst_mult_4_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_152 (
// Equation(s):
// Xd_0__inst_mult_5_520  = SUM(( GND ) + ( Xd_0__inst_mult_5_506  ) + ( Xd_0__inst_mult_5_505  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_505 ),
	.sharein(Xd_0__inst_mult_5_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_520 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_153 (
// Equation(s):
// Xd_0__inst_mult_5_524  = SUM(( (din_a[69] & din_b[65]) ) + ( Xd_0__inst_mult_5_510  ) + ( Xd_0__inst_mult_5_509  ))
// Xd_0__inst_mult_5_525  = CARRY(( (din_a[69] & din_b[65]) ) + ( Xd_0__inst_mult_5_510  ) + ( Xd_0__inst_mult_5_509  ))
// Xd_0__inst_mult_5_526  = SHARE((din_a[69] & din_b[66]))

	.dataa(!din_a[69]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_509 ),
	.sharein(Xd_0__inst_mult_5_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_524 ),
	.cout(Xd_0__inst_mult_5_525 ),
	.shareout(Xd_0__inst_mult_5_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_154 (
// Equation(s):
// Xd_0__inst_mult_5_528  = SUM(( (din_a[65] & din_b[69]) ) + ( Xd_0__inst_mult_5_514  ) + ( Xd_0__inst_mult_5_513  ))
// Xd_0__inst_mult_5_529  = CARRY(( (din_a[65] & din_b[69]) ) + ( Xd_0__inst_mult_5_514  ) + ( Xd_0__inst_mult_5_513  ))
// Xd_0__inst_mult_5_530  = SHARE((din_a[65] & din_b[70]))

	.dataa(!din_a[65]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_513 ),
	.sharein(Xd_0__inst_mult_5_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_528 ),
	.cout(Xd_0__inst_mult_5_529 ),
	.shareout(Xd_0__inst_mult_5_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_155 (
// Equation(s):
// Xd_0__inst_mult_5_532  = SUM(( (!din_a[67] & (((din_a[66] & din_b[68])))) # (din_a[67] & (!din_b[67] $ (((!din_a[66]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_518  ) + ( Xd_0__inst_mult_5_517  ))
// Xd_0__inst_mult_5_533  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[68])))) # (din_a[67] & (!din_b[67] $ (((!din_a[66]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_518  ) + ( Xd_0__inst_mult_5_517  ))
// Xd_0__inst_mult_5_534  = SHARE((din_a[67] & (din_b[67] & (din_a[66] & din_b[68]))))

	.dataa(!din_a[67]),
	.datab(!din_b[67]),
	.datac(!din_a[66]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_517 ),
	.sharein(Xd_0__inst_mult_5_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_532 ),
	.cout(Xd_0__inst_mult_5_533 ),
	.shareout(Xd_0__inst_mult_5_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_156 (
// Equation(s):
// Xd_0__inst_mult_2_524  = SUM(( GND ) + ( Xd_0__inst_mult_2_510  ) + ( Xd_0__inst_mult_2_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_509 ),
	.sharein(Xd_0__inst_mult_2_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_524 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_157 (
// Equation(s):
// Xd_0__inst_mult_2_528  = SUM(( (din_a[33] & din_b[29]) ) + ( Xd_0__inst_mult_2_514  ) + ( Xd_0__inst_mult_2_513  ))
// Xd_0__inst_mult_2_529  = CARRY(( (din_a[33] & din_b[29]) ) + ( Xd_0__inst_mult_2_514  ) + ( Xd_0__inst_mult_2_513  ))
// Xd_0__inst_mult_2_530  = SHARE((din_a[33] & din_b[30]))

	.dataa(!din_a[33]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_513 ),
	.sharein(Xd_0__inst_mult_2_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_528 ),
	.cout(Xd_0__inst_mult_2_529 ),
	.shareout(Xd_0__inst_mult_2_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_158 (
// Equation(s):
// Xd_0__inst_mult_2_532  = SUM(( (din_a[29] & din_b[33]) ) + ( Xd_0__inst_mult_2_518  ) + ( Xd_0__inst_mult_2_517  ))
// Xd_0__inst_mult_2_533  = CARRY(( (din_a[29] & din_b[33]) ) + ( Xd_0__inst_mult_2_518  ) + ( Xd_0__inst_mult_2_517  ))
// Xd_0__inst_mult_2_534  = SHARE((din_a[29] & din_b[34]))

	.dataa(!din_a[29]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_517 ),
	.sharein(Xd_0__inst_mult_2_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_532 ),
	.cout(Xd_0__inst_mult_2_533 ),
	.shareout(Xd_0__inst_mult_2_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_159 (
// Equation(s):
// Xd_0__inst_mult_2_536  = SUM(( (!din_a[31] & (((din_a[30] & din_b[32])))) # (din_a[31] & (!din_b[31] $ (((!din_a[30]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_522  ) + ( Xd_0__inst_mult_2_521  ))
// Xd_0__inst_mult_2_537  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[32])))) # (din_a[31] & (!din_b[31] $ (((!din_a[30]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_522  ) + ( Xd_0__inst_mult_2_521  ))
// Xd_0__inst_mult_2_538  = SHARE((din_a[31] & (din_b[31] & (din_a[30] & din_b[32]))))

	.dataa(!din_a[31]),
	.datab(!din_b[31]),
	.datac(!din_a[30]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_521 ),
	.sharein(Xd_0__inst_mult_2_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_536 ),
	.cout(Xd_0__inst_mult_2_537 ),
	.shareout(Xd_0__inst_mult_2_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_152 (
// Equation(s):
// Xd_0__inst_mult_3_520  = SUM(( GND ) + ( Xd_0__inst_mult_3_506  ) + ( Xd_0__inst_mult_3_505  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_505 ),
	.sharein(Xd_0__inst_mult_3_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_520 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_153 (
// Equation(s):
// Xd_0__inst_mult_3_524  = SUM(( (din_a[45] & din_b[41]) ) + ( Xd_0__inst_mult_3_510  ) + ( Xd_0__inst_mult_3_509  ))
// Xd_0__inst_mult_3_525  = CARRY(( (din_a[45] & din_b[41]) ) + ( Xd_0__inst_mult_3_510  ) + ( Xd_0__inst_mult_3_509  ))
// Xd_0__inst_mult_3_526  = SHARE((din_a[45] & din_b[42]))

	.dataa(!din_a[45]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_509 ),
	.sharein(Xd_0__inst_mult_3_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_524 ),
	.cout(Xd_0__inst_mult_3_525 ),
	.shareout(Xd_0__inst_mult_3_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_154 (
// Equation(s):
// Xd_0__inst_mult_3_528  = SUM(( (din_a[41] & din_b[45]) ) + ( Xd_0__inst_mult_3_514  ) + ( Xd_0__inst_mult_3_513  ))
// Xd_0__inst_mult_3_529  = CARRY(( (din_a[41] & din_b[45]) ) + ( Xd_0__inst_mult_3_514  ) + ( Xd_0__inst_mult_3_513  ))
// Xd_0__inst_mult_3_530  = SHARE((din_a[41] & din_b[46]))

	.dataa(!din_a[41]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_513 ),
	.sharein(Xd_0__inst_mult_3_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_528 ),
	.cout(Xd_0__inst_mult_3_529 ),
	.shareout(Xd_0__inst_mult_3_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_155 (
// Equation(s):
// Xd_0__inst_mult_3_532  = SUM(( (!din_a[43] & (((din_a[42] & din_b[44])))) # (din_a[43] & (!din_b[43] $ (((!din_a[42]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_518  ) + ( Xd_0__inst_mult_3_517  ))
// Xd_0__inst_mult_3_533  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[44])))) # (din_a[43] & (!din_b[43] $ (((!din_a[42]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_518  ) + ( Xd_0__inst_mult_3_517  ))
// Xd_0__inst_mult_3_534  = SHARE((din_a[43] & (din_b[43] & (din_a[42] & din_b[44]))))

	.dataa(!din_a[43]),
	.datab(!din_b[43]),
	.datac(!din_a[42]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_517 ),
	.sharein(Xd_0__inst_mult_3_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_532 ),
	.cout(Xd_0__inst_mult_3_533 ),
	.shareout(Xd_0__inst_mult_3_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_156 (
// Equation(s):
// Xd_0__inst_mult_0_524  = SUM(( GND ) + ( Xd_0__inst_mult_0_510  ) + ( Xd_0__inst_mult_0_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_509 ),
	.sharein(Xd_0__inst_mult_0_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_524 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_157 (
// Equation(s):
// Xd_0__inst_mult_0_528  = SUM(( (din_a[9] & din_b[5]) ) + ( Xd_0__inst_mult_0_514  ) + ( Xd_0__inst_mult_0_513  ))
// Xd_0__inst_mult_0_529  = CARRY(( (din_a[9] & din_b[5]) ) + ( Xd_0__inst_mult_0_514  ) + ( Xd_0__inst_mult_0_513  ))
// Xd_0__inst_mult_0_530  = SHARE((din_a[9] & din_b[6]))

	.dataa(!din_a[9]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_513 ),
	.sharein(Xd_0__inst_mult_0_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_528 ),
	.cout(Xd_0__inst_mult_0_529 ),
	.shareout(Xd_0__inst_mult_0_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_158 (
// Equation(s):
// Xd_0__inst_mult_0_532  = SUM(( (din_a[5] & din_b[9]) ) + ( Xd_0__inst_mult_0_518  ) + ( Xd_0__inst_mult_0_517  ))
// Xd_0__inst_mult_0_533  = CARRY(( (din_a[5] & din_b[9]) ) + ( Xd_0__inst_mult_0_518  ) + ( Xd_0__inst_mult_0_517  ))
// Xd_0__inst_mult_0_534  = SHARE((din_a[5] & din_b[10]))

	.dataa(!din_a[5]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_517 ),
	.sharein(Xd_0__inst_mult_0_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_532 ),
	.cout(Xd_0__inst_mult_0_533 ),
	.shareout(Xd_0__inst_mult_0_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_159 (
// Equation(s):
// Xd_0__inst_mult_0_536  = SUM(( (!din_a[7] & (((din_a[6] & din_b[8])))) # (din_a[7] & (!din_b[7] $ (((!din_a[6]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_522  ) + ( Xd_0__inst_mult_0_521  ))
// Xd_0__inst_mult_0_537  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[8])))) # (din_a[7] & (!din_b[7] $ (((!din_a[6]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_522  ) + ( Xd_0__inst_mult_0_521  ))
// Xd_0__inst_mult_0_538  = SHARE((din_a[7] & (din_b[7] & (din_a[6] & din_b[8]))))

	.dataa(!din_a[7]),
	.datab(!din_b[7]),
	.datac(!din_a[6]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_521 ),
	.sharein(Xd_0__inst_mult_0_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_536 ),
	.cout(Xd_0__inst_mult_0_537 ),
	.shareout(Xd_0__inst_mult_0_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_156 (
// Equation(s):
// Xd_0__inst_mult_1_524  = SUM(( GND ) + ( Xd_0__inst_mult_1_510  ) + ( Xd_0__inst_mult_1_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_509 ),
	.sharein(Xd_0__inst_mult_1_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_524 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_157 (
// Equation(s):
// Xd_0__inst_mult_1_528  = SUM(( (din_a[21] & din_b[17]) ) + ( Xd_0__inst_mult_1_514  ) + ( Xd_0__inst_mult_1_513  ))
// Xd_0__inst_mult_1_529  = CARRY(( (din_a[21] & din_b[17]) ) + ( Xd_0__inst_mult_1_514  ) + ( Xd_0__inst_mult_1_513  ))
// Xd_0__inst_mult_1_530  = SHARE((din_a[21] & din_b[18]))

	.dataa(!din_a[21]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_513 ),
	.sharein(Xd_0__inst_mult_1_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_528 ),
	.cout(Xd_0__inst_mult_1_529 ),
	.shareout(Xd_0__inst_mult_1_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_158 (
// Equation(s):
// Xd_0__inst_mult_1_532  = SUM(( (din_a[17] & din_b[21]) ) + ( Xd_0__inst_mult_1_518  ) + ( Xd_0__inst_mult_1_517  ))
// Xd_0__inst_mult_1_533  = CARRY(( (din_a[17] & din_b[21]) ) + ( Xd_0__inst_mult_1_518  ) + ( Xd_0__inst_mult_1_517  ))
// Xd_0__inst_mult_1_534  = SHARE((din_a[17] & din_b[22]))

	.dataa(!din_a[17]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_517 ),
	.sharein(Xd_0__inst_mult_1_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_532 ),
	.cout(Xd_0__inst_mult_1_533 ),
	.shareout(Xd_0__inst_mult_1_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_159 (
// Equation(s):
// Xd_0__inst_mult_1_536  = SUM(( (!din_a[19] & (((din_a[18] & din_b[20])))) # (din_a[19] & (!din_b[19] $ (((!din_a[18]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_522  ) + ( Xd_0__inst_mult_1_521  ))
// Xd_0__inst_mult_1_537  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[20])))) # (din_a[19] & (!din_b[19] $ (((!din_a[18]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_522  ) + ( Xd_0__inst_mult_1_521  ))
// Xd_0__inst_mult_1_538  = SHARE((din_a[19] & (din_b[19] & (din_a[18] & din_b[20]))))

	.dataa(!din_a[19]),
	.datab(!din_b[19]),
	.datac(!din_a[18]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_521 ),
	.sharein(Xd_0__inst_mult_1_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_536 ),
	.cout(Xd_0__inst_mult_1_537 ),
	.shareout(Xd_0__inst_mult_1_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_161 (
// Equation(s):
// Xd_0__inst_mult_12_556  = SUM(( (din_a[152] & din_b[151]) ) + ( Xd_0__inst_mult_12_550  ) + ( Xd_0__inst_mult_12_549  ))
// Xd_0__inst_mult_12_557  = CARRY(( (din_a[152] & din_b[151]) ) + ( Xd_0__inst_mult_12_550  ) + ( Xd_0__inst_mult_12_549  ))
// Xd_0__inst_mult_12_558  = SHARE((din_b[151] & din_a[153]))

	.dataa(!din_a[152]),
	.datab(!din_b[151]),
	.datac(!din_a[153]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_549 ),
	.sharein(Xd_0__inst_mult_12_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_556 ),
	.cout(Xd_0__inst_mult_12_557 ),
	.shareout(Xd_0__inst_mult_12_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_160 (
// Equation(s):
// Xd_0__inst_mult_14_540  = SUM(( GND ) + ( Xd_0__inst_mult_12_554  ) + ( Xd_0__inst_mult_12_553  ))
// Xd_0__inst_mult_14_541  = CARRY(( GND ) + ( Xd_0__inst_mult_12_554  ) + ( Xd_0__inst_mult_12_553  ))
// Xd_0__inst_mult_14_542  = SHARE(VCC)

	.dataa(!din_a[170]),
	.datab(!din_b[175]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_553 ),
	.sharein(Xd_0__inst_mult_12_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_540 ),
	.cout(Xd_0__inst_mult_14_541 ),
	.shareout(Xd_0__inst_mult_14_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_160 (
// Equation(s):
// Xd_0__inst_mult_13_540  = SUM(( (din_a[164] & din_b[163]) ) + ( Xd_0__inst_mult_13_530  ) + ( Xd_0__inst_mult_13_529  ))
// Xd_0__inst_mult_13_541  = CARRY(( (din_a[164] & din_b[163]) ) + ( Xd_0__inst_mult_13_530  ) + ( Xd_0__inst_mult_13_529  ))
// Xd_0__inst_mult_13_542  = SHARE((din_b[163] & din_a[165]))

	.dataa(!din_a[164]),
	.datab(!din_b[163]),
	.datac(!din_a[165]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_529 ),
	.sharein(Xd_0__inst_mult_13_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_540 ),
	.cout(Xd_0__inst_mult_13_541 ),
	.shareout(Xd_0__inst_mult_13_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_161 (
// Equation(s):
// Xd_0__inst_mult_13_544  = SUM(( (!din_a[163] & (((din_a[162] & din_b[165])))) # (din_a[163] & (!din_b[164] $ (((!din_a[162]) # (!din_b[165]))))) ) + ( Xd_0__inst_mult_13_534  ) + ( Xd_0__inst_mult_13_533  ))
// Xd_0__inst_mult_13_545  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[165])))) # (din_a[163] & (!din_b[164] $ (((!din_a[162]) # (!din_b[165]))))) ) + ( Xd_0__inst_mult_13_534  ) + ( Xd_0__inst_mult_13_533  ))
// Xd_0__inst_mult_13_546  = SHARE((din_a[163] & (din_b[164] & (din_a[162] & din_b[165]))))

	.dataa(!din_a[163]),
	.datab(!din_b[164]),
	.datac(!din_a[162]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_533 ),
	.sharein(Xd_0__inst_mult_13_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_544 ),
	.cout(Xd_0__inst_mult_13_545 ),
	.shareout(Xd_0__inst_mult_13_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_160 (
// Equation(s):
// Xd_0__inst_mult_1_540  = SUM(( GND ) + ( Xd_0__inst_mult_13_538  ) + ( Xd_0__inst_mult_13_537  ))
// Xd_0__inst_mult_1_541  = CARRY(( GND ) + ( Xd_0__inst_mult_13_538  ) + ( Xd_0__inst_mult_13_537  ))
// Xd_0__inst_mult_1_542  = SHARE(VCC)

	.dataa(!din_a[15]),
	.datab(!din_b[13]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_537 ),
	.sharein(Xd_0__inst_mult_13_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_540 ),
	.cout(Xd_0__inst_mult_1_541 ),
	.shareout(Xd_0__inst_mult_1_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_161 (
// Equation(s):
// Xd_0__inst_mult_14_544  = SUM(( (din_a[176] & din_b[175]) ) + ( Xd_0__inst_mult_14_530  ) + ( Xd_0__inst_mult_14_529  ))
// Xd_0__inst_mult_14_545  = CARRY(( (din_a[176] & din_b[175]) ) + ( Xd_0__inst_mult_14_530  ) + ( Xd_0__inst_mult_14_529  ))
// Xd_0__inst_mult_14_546  = SHARE((din_b[175] & din_a[177]))

	.dataa(!din_a[176]),
	.datab(!din_b[175]),
	.datac(!din_a[177]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_529 ),
	.sharein(Xd_0__inst_mult_14_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_544 ),
	.cout(Xd_0__inst_mult_14_545 ),
	.shareout(Xd_0__inst_mult_14_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_162 (
// Equation(s):
// Xd_0__inst_mult_14_548  = SUM(( (!din_a[175] & (((din_a[174] & din_b[177])))) # (din_a[175] & (!din_b[176] $ (((!din_a[174]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_14_534  ) + ( Xd_0__inst_mult_14_533  ))
// Xd_0__inst_mult_14_549  = CARRY(( (!din_a[175] & (((din_a[174] & din_b[177])))) # (din_a[175] & (!din_b[176] $ (((!din_a[174]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_14_534  ) + ( Xd_0__inst_mult_14_533  ))
// Xd_0__inst_mult_14_550  = SHARE((din_a[175] & (din_b[176] & (din_a[174] & din_b[177]))))

	.dataa(!din_a[175]),
	.datab(!din_b[176]),
	.datac(!din_a[174]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_533 ),
	.sharein(Xd_0__inst_mult_14_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_548 ),
	.cout(Xd_0__inst_mult_14_549 ),
	.shareout(Xd_0__inst_mult_14_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_165 (
// Equation(s):
// Xd_0__inst_mult_15_560  = SUM(( GND ) + ( Xd_0__inst_mult_14_538  ) + ( Xd_0__inst_mult_14_537  ))
// Xd_0__inst_mult_15_561  = CARRY(( GND ) + ( Xd_0__inst_mult_14_538  ) + ( Xd_0__inst_mult_14_537  ))
// Xd_0__inst_mult_15_562  = SHARE(VCC)

	.dataa(!din_a[183]),
	.datab(!din_b[181]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_537 ),
	.sharein(Xd_0__inst_mult_14_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_560 ),
	.cout(Xd_0__inst_mult_15_561 ),
	.shareout(Xd_0__inst_mult_15_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_166 (
// Equation(s):
// Xd_0__inst_mult_15_564  = SUM(( (din_a[188] & din_b[187]) ) + ( Xd_0__inst_mult_15_554  ) + ( Xd_0__inst_mult_15_553  ))
// Xd_0__inst_mult_15_565  = CARRY(( (din_a[188] & din_b[187]) ) + ( Xd_0__inst_mult_15_554  ) + ( Xd_0__inst_mult_15_553  ))
// Xd_0__inst_mult_15_566  = SHARE((din_b[187] & din_a[189]))

	.dataa(!din_a[188]),
	.datab(!din_b[187]),
	.datac(!din_a[189]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_553 ),
	.sharein(Xd_0__inst_mult_15_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_564 ),
	.cout(Xd_0__inst_mult_15_565 ),
	.shareout(Xd_0__inst_mult_15_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_163 (
// Equation(s):
// Xd_0__inst_mult_14_552  = SUM(( GND ) + ( Xd_0__inst_mult_15_558  ) + ( Xd_0__inst_mult_15_557  ))
// Xd_0__inst_mult_14_553  = CARRY(( GND ) + ( Xd_0__inst_mult_15_558  ) + ( Xd_0__inst_mult_15_557  ))
// Xd_0__inst_mult_14_554  = SHARE(VCC)

	.dataa(!din_a[171]),
	.datab(!din_b[169]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_557 ),
	.sharein(Xd_0__inst_mult_15_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_552 ),
	.cout(Xd_0__inst_mult_14_553 ),
	.shareout(Xd_0__inst_mult_14_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_156 (
// Equation(s):
// Xd_0__inst_mult_10_536  = SUM(( (din_a[128] & din_b[127]) ) + ( Xd_0__inst_mult_10_526  ) + ( Xd_0__inst_mult_10_525  ))
// Xd_0__inst_mult_10_537  = CARRY(( (din_a[128] & din_b[127]) ) + ( Xd_0__inst_mult_10_526  ) + ( Xd_0__inst_mult_10_525  ))
// Xd_0__inst_mult_10_538  = SHARE((din_b[127] & din_a[129]))

	.dataa(!din_a[128]),
	.datab(!din_b[127]),
	.datac(!din_a[129]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_525 ),
	.sharein(Xd_0__inst_mult_10_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_536 ),
	.cout(Xd_0__inst_mult_10_537 ),
	.shareout(Xd_0__inst_mult_10_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_157 (
// Equation(s):
// Xd_0__inst_mult_10_540  = SUM(( (!din_a[127] & (((din_a[126] & din_b[129])))) # (din_a[127] & (!din_b[128] $ (((!din_a[126]) # (!din_b[129]))))) ) + ( Xd_0__inst_mult_10_530  ) + ( Xd_0__inst_mult_10_529  ))
// Xd_0__inst_mult_10_541  = CARRY(( (!din_a[127] & (((din_a[126] & din_b[129])))) # (din_a[127] & (!din_b[128] $ (((!din_a[126]) # (!din_b[129]))))) ) + ( Xd_0__inst_mult_10_530  ) + ( Xd_0__inst_mult_10_529  ))
// Xd_0__inst_mult_10_542  = SHARE((din_a[127] & (din_b[128] & (din_a[126] & din_b[129]))))

	.dataa(!din_a[127]),
	.datab(!din_b[128]),
	.datac(!din_a[126]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_529 ),
	.sharein(Xd_0__inst_mult_10_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_540 ),
	.cout(Xd_0__inst_mult_10_541 ),
	.shareout(Xd_0__inst_mult_10_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_160 (
// Equation(s):
// Xd_0__inst_mult_0_540  = SUM(( GND ) + ( Xd_0__inst_mult_10_534  ) + ( Xd_0__inst_mult_10_533  ))
// Xd_0__inst_mult_0_541  = CARRY(( GND ) + ( Xd_0__inst_mult_10_534  ) + ( Xd_0__inst_mult_10_533  ))
// Xd_0__inst_mult_0_542  = SHARE(VCC)

	.dataa(!din_a[2]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_533 ),
	.sharein(Xd_0__inst_mult_10_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_540 ),
	.cout(Xd_0__inst_mult_0_541 ),
	.shareout(Xd_0__inst_mult_0_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_160 (
// Equation(s):
// Xd_0__inst_mult_11_540  = SUM(( (din_a[140] & din_b[139]) ) + ( Xd_0__inst_mult_11_530  ) + ( Xd_0__inst_mult_11_529  ))
// Xd_0__inst_mult_11_541  = CARRY(( (din_a[140] & din_b[139]) ) + ( Xd_0__inst_mult_11_530  ) + ( Xd_0__inst_mult_11_529  ))
// Xd_0__inst_mult_11_542  = SHARE((din_b[139] & din_a[141]))

	.dataa(!din_a[140]),
	.datab(!din_b[139]),
	.datac(!din_a[141]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_529 ),
	.sharein(Xd_0__inst_mult_11_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_540 ),
	.cout(Xd_0__inst_mult_11_541 ),
	.shareout(Xd_0__inst_mult_11_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_161 (
// Equation(s):
// Xd_0__inst_mult_11_544  = SUM(( (!din_a[139] & (((din_a[138] & din_b[141])))) # (din_a[139] & (!din_b[140] $ (((!din_a[138]) # (!din_b[141]))))) ) + ( Xd_0__inst_mult_11_534  ) + ( Xd_0__inst_mult_11_533  ))
// Xd_0__inst_mult_11_545  = CARRY(( (!din_a[139] & (((din_a[138] & din_b[141])))) # (din_a[139] & (!din_b[140] $ (((!din_a[138]) # (!din_b[141]))))) ) + ( Xd_0__inst_mult_11_534  ) + ( Xd_0__inst_mult_11_533  ))
// Xd_0__inst_mult_11_546  = SHARE((din_a[139] & (din_b[140] & (din_a[138] & din_b[141]))))

	.dataa(!din_a[139]),
	.datab(!din_b[140]),
	.datac(!din_a[138]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_533 ),
	.sharein(Xd_0__inst_mult_11_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_544 ),
	.cout(Xd_0__inst_mult_11_545 ),
	.shareout(Xd_0__inst_mult_11_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_156 (
// Equation(s):
// Xd_0__inst_mult_3_536  = SUM(( GND ) + ( Xd_0__inst_mult_11_538  ) + ( Xd_0__inst_mult_11_537  ))
// Xd_0__inst_mult_3_537  = CARRY(( GND ) + ( Xd_0__inst_mult_11_538  ) + ( Xd_0__inst_mult_11_537  ))
// Xd_0__inst_mult_3_538  = SHARE(VCC)

	.dataa(!din_a[38]),
	.datab(!din_b[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_537 ),
	.sharein(Xd_0__inst_mult_11_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_536 ),
	.cout(Xd_0__inst_mult_3_537 ),
	.shareout(Xd_0__inst_mult_3_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_160 (
// Equation(s):
// Xd_0__inst_mult_8_540  = SUM(( (din_a[104] & din_b[103]) ) + ( Xd_0__inst_mult_8_530  ) + ( Xd_0__inst_mult_8_529  ))
// Xd_0__inst_mult_8_541  = CARRY(( (din_a[104] & din_b[103]) ) + ( Xd_0__inst_mult_8_530  ) + ( Xd_0__inst_mult_8_529  ))
// Xd_0__inst_mult_8_542  = SHARE((din_b[103] & din_a[105]))

	.dataa(!din_a[104]),
	.datab(!din_b[103]),
	.datac(!din_a[105]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_529 ),
	.sharein(Xd_0__inst_mult_8_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_540 ),
	.cout(Xd_0__inst_mult_8_541 ),
	.shareout(Xd_0__inst_mult_8_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_161 (
// Equation(s):
// Xd_0__inst_mult_8_544  = SUM(( (!din_a[103] & (((din_a[102] & din_b[105])))) # (din_a[103] & (!din_b[104] $ (((!din_a[102]) # (!din_b[105]))))) ) + ( Xd_0__inst_mult_8_534  ) + ( Xd_0__inst_mult_8_533  ))
// Xd_0__inst_mult_8_545  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[105])))) # (din_a[103] & (!din_b[104] $ (((!din_a[102]) # (!din_b[105]))))) ) + ( Xd_0__inst_mult_8_534  ) + ( Xd_0__inst_mult_8_533  ))
// Xd_0__inst_mult_8_546  = SHARE((din_a[103] & (din_b[104] & (din_a[102] & din_b[105]))))

	.dataa(!din_a[103]),
	.datab(!din_b[104]),
	.datac(!din_a[102]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_533 ),
	.sharein(Xd_0__inst_mult_8_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_544 ),
	.cout(Xd_0__inst_mult_8_545 ),
	.shareout(Xd_0__inst_mult_8_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_160 (
// Equation(s):
// Xd_0__inst_mult_2_540  = SUM(( GND ) + ( Xd_0__inst_mult_8_538  ) + ( Xd_0__inst_mult_8_537  ))
// Xd_0__inst_mult_2_541  = CARRY(( GND ) + ( Xd_0__inst_mult_8_538  ) + ( Xd_0__inst_mult_8_537  ))
// Xd_0__inst_mult_2_542  = SHARE(VCC)

	.dataa(!din_a[26]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_537 ),
	.sharein(Xd_0__inst_mult_8_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_540 ),
	.cout(Xd_0__inst_mult_2_541 ),
	.shareout(Xd_0__inst_mult_2_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_156 (
// Equation(s):
// Xd_0__inst_mult_9_536  = SUM(( (din_a[116] & din_b[115]) ) + ( Xd_0__inst_mult_9_526  ) + ( Xd_0__inst_mult_9_525  ))
// Xd_0__inst_mult_9_537  = CARRY(( (din_a[116] & din_b[115]) ) + ( Xd_0__inst_mult_9_526  ) + ( Xd_0__inst_mult_9_525  ))
// Xd_0__inst_mult_9_538  = SHARE((din_b[115] & din_a[117]))

	.dataa(!din_a[116]),
	.datab(!din_b[115]),
	.datac(!din_a[117]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_525 ),
	.sharein(Xd_0__inst_mult_9_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_536 ),
	.cout(Xd_0__inst_mult_9_537 ),
	.shareout(Xd_0__inst_mult_9_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_157 (
// Equation(s):
// Xd_0__inst_mult_9_540  = SUM(( (!din_a[115] & (((din_a[114] & din_b[117])))) # (din_a[115] & (!din_b[116] $ (((!din_a[114]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_9_530  ) + ( Xd_0__inst_mult_9_529  ))
// Xd_0__inst_mult_9_541  = CARRY(( (!din_a[115] & (((din_a[114] & din_b[117])))) # (din_a[115] & (!din_b[116] $ (((!din_a[114]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_9_530  ) + ( Xd_0__inst_mult_9_529  ))
// Xd_0__inst_mult_9_542  = SHARE((din_a[115] & (din_b[116] & (din_a[114] & din_b[117]))))

	.dataa(!din_a[115]),
	.datab(!din_b[116]),
	.datac(!din_a[114]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_529 ),
	.sharein(Xd_0__inst_mult_9_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_540 ),
	.cout(Xd_0__inst_mult_9_541 ),
	.shareout(Xd_0__inst_mult_9_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_161 (
// Equation(s):
// Xd_0__inst_mult_1_544  = SUM(( GND ) + ( Xd_0__inst_mult_9_534  ) + ( Xd_0__inst_mult_9_533  ))
// Xd_0__inst_mult_1_545  = CARRY(( GND ) + ( Xd_0__inst_mult_9_534  ) + ( Xd_0__inst_mult_9_533  ))
// Xd_0__inst_mult_1_546  = SHARE(VCC)

	.dataa(!din_a[14]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_533 ),
	.sharein(Xd_0__inst_mult_9_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_544 ),
	.cout(Xd_0__inst_mult_1_545 ),
	.shareout(Xd_0__inst_mult_1_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_156 (
// Equation(s):
// Xd_0__inst_mult_6_536  = SUM(( (din_a[80] & din_b[79]) ) + ( Xd_0__inst_mult_6_526  ) + ( Xd_0__inst_mult_6_525  ))
// Xd_0__inst_mult_6_537  = CARRY(( (din_a[80] & din_b[79]) ) + ( Xd_0__inst_mult_6_526  ) + ( Xd_0__inst_mult_6_525  ))
// Xd_0__inst_mult_6_538  = SHARE((din_b[79] & din_a[81]))

	.dataa(!din_a[80]),
	.datab(!din_b[79]),
	.datac(!din_a[81]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_525 ),
	.sharein(Xd_0__inst_mult_6_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_536 ),
	.cout(Xd_0__inst_mult_6_537 ),
	.shareout(Xd_0__inst_mult_6_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_157 (
// Equation(s):
// Xd_0__inst_mult_6_540  = SUM(( (!din_a[79] & (((din_a[78] & din_b[81])))) # (din_a[79] & (!din_b[80] $ (((!din_a[78]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_6_530  ) + ( Xd_0__inst_mult_6_529  ))
// Xd_0__inst_mult_6_541  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[81])))) # (din_a[79] & (!din_b[80] $ (((!din_a[78]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_6_530  ) + ( Xd_0__inst_mult_6_529  ))
// Xd_0__inst_mult_6_542  = SHARE((din_a[79] & (din_b[80] & (din_a[78] & din_b[81]))))

	.dataa(!din_a[79]),
	.datab(!din_b[80]),
	.datac(!din_a[78]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_529 ),
	.sharein(Xd_0__inst_mult_6_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_540 ),
	.cout(Xd_0__inst_mult_6_541 ),
	.shareout(Xd_0__inst_mult_6_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_156 (
// Equation(s):
// Xd_0__inst_mult_5_536  = SUM(( GND ) + ( Xd_0__inst_mult_6_534  ) + ( Xd_0__inst_mult_6_533  ))
// Xd_0__inst_mult_5_537  = CARRY(( GND ) + ( Xd_0__inst_mult_6_534  ) + ( Xd_0__inst_mult_6_533  ))
// Xd_0__inst_mult_5_538  = SHARE(VCC)

	.dataa(!din_a[62]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_533 ),
	.sharein(Xd_0__inst_mult_6_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_536 ),
	.cout(Xd_0__inst_mult_5_537 ),
	.shareout(Xd_0__inst_mult_5_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_156 (
// Equation(s):
// Xd_0__inst_mult_7_536  = SUM(( (din_a[92] & din_b[91]) ) + ( Xd_0__inst_mult_7_526  ) + ( Xd_0__inst_mult_7_525  ))
// Xd_0__inst_mult_7_537  = CARRY(( (din_a[92] & din_b[91]) ) + ( Xd_0__inst_mult_7_526  ) + ( Xd_0__inst_mult_7_525  ))
// Xd_0__inst_mult_7_538  = SHARE((din_b[91] & din_a[93]))

	.dataa(!din_a[92]),
	.datab(!din_b[91]),
	.datac(!din_a[93]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_525 ),
	.sharein(Xd_0__inst_mult_7_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_536 ),
	.cout(Xd_0__inst_mult_7_537 ),
	.shareout(Xd_0__inst_mult_7_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_157 (
// Equation(s):
// Xd_0__inst_mult_7_540  = SUM(( (!din_a[91] & (((din_a[90] & din_b[93])))) # (din_a[91] & (!din_b[92] $ (((!din_a[90]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_7_530  ) + ( Xd_0__inst_mult_7_529  ))
// Xd_0__inst_mult_7_541  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[93])))) # (din_a[91] & (!din_b[92] $ (((!din_a[90]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_7_530  ) + ( Xd_0__inst_mult_7_529  ))
// Xd_0__inst_mult_7_542  = SHARE((din_a[91] & (din_b[92] & (din_a[90] & din_b[93]))))

	.dataa(!din_a[91]),
	.datab(!din_b[92]),
	.datac(!din_a[90]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_529 ),
	.sharein(Xd_0__inst_mult_7_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_540 ),
	.cout(Xd_0__inst_mult_7_541 ),
	.shareout(Xd_0__inst_mult_7_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_158 (
// Equation(s):
// Xd_0__inst_mult_7_544  = SUM(( GND ) + ( Xd_0__inst_mult_7_534  ) + ( Xd_0__inst_mult_7_533  ))
// Xd_0__inst_mult_7_545  = CARRY(( GND ) + ( Xd_0__inst_mult_7_534  ) + ( Xd_0__inst_mult_7_533  ))
// Xd_0__inst_mult_7_546  = SHARE(VCC)

	.dataa(!din_a[86]),
	.datab(!din_b[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_533 ),
	.sharein(Xd_0__inst_mult_7_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_544 ),
	.cout(Xd_0__inst_mult_7_545 ),
	.shareout(Xd_0__inst_mult_7_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_165 (
// Equation(s):
// Xd_0__inst_mult_4_560  = SUM(( (din_a[56] & din_b[55]) ) + ( Xd_0__inst_mult_4_554  ) + ( Xd_0__inst_mult_4_553  ))
// Xd_0__inst_mult_4_561  = CARRY(( (din_a[56] & din_b[55]) ) + ( Xd_0__inst_mult_4_554  ) + ( Xd_0__inst_mult_4_553  ))
// Xd_0__inst_mult_4_562  = SHARE((din_b[55] & din_a[57]))

	.dataa(!din_a[56]),
	.datab(!din_b[55]),
	.datac(!din_a[57]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_553 ),
	.sharein(Xd_0__inst_mult_4_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_560 ),
	.cout(Xd_0__inst_mult_4_561 ),
	.shareout(Xd_0__inst_mult_4_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_158 (
// Equation(s):
// Xd_0__inst_mult_6_544  = SUM(( GND ) + ( Xd_0__inst_mult_4_558  ) + ( Xd_0__inst_mult_4_557  ))
// Xd_0__inst_mult_6_545  = CARRY(( GND ) + ( Xd_0__inst_mult_4_558  ) + ( Xd_0__inst_mult_4_557  ))
// Xd_0__inst_mult_6_546  = SHARE(VCC)

	.dataa(!din_a[74]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_557 ),
	.sharein(Xd_0__inst_mult_4_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_544 ),
	.cout(Xd_0__inst_mult_6_545 ),
	.shareout(Xd_0__inst_mult_6_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_157 (
// Equation(s):
// Xd_0__inst_mult_5_540  = SUM(( (din_a[68] & din_b[67]) ) + ( Xd_0__inst_mult_5_526  ) + ( Xd_0__inst_mult_5_525  ))
// Xd_0__inst_mult_5_541  = CARRY(( (din_a[68] & din_b[67]) ) + ( Xd_0__inst_mult_5_526  ) + ( Xd_0__inst_mult_5_525  ))
// Xd_0__inst_mult_5_542  = SHARE((din_b[67] & din_a[69]))

	.dataa(!din_a[68]),
	.datab(!din_b[67]),
	.datac(!din_a[69]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_525 ),
	.sharein(Xd_0__inst_mult_5_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_540 ),
	.cout(Xd_0__inst_mult_5_541 ),
	.shareout(Xd_0__inst_mult_5_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_158 (
// Equation(s):
// Xd_0__inst_mult_5_544  = SUM(( (!din_a[67] & (((din_a[66] & din_b[69])))) # (din_a[67] & (!din_b[68] $ (((!din_a[66]) # (!din_b[69]))))) ) + ( Xd_0__inst_mult_5_530  ) + ( Xd_0__inst_mult_5_529  ))
// Xd_0__inst_mult_5_545  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[69])))) # (din_a[67] & (!din_b[68] $ (((!din_a[66]) # (!din_b[69]))))) ) + ( Xd_0__inst_mult_5_530  ) + ( Xd_0__inst_mult_5_529  ))
// Xd_0__inst_mult_5_546  = SHARE((din_a[67] & (din_b[68] & (din_a[66] & din_b[69]))))

	.dataa(!din_a[67]),
	.datab(!din_b[68]),
	.datac(!din_a[66]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_529 ),
	.sharein(Xd_0__inst_mult_5_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_544 ),
	.cout(Xd_0__inst_mult_5_545 ),
	.shareout(Xd_0__inst_mult_5_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_158 (
// Equation(s):
// Xd_0__inst_mult_9_544  = SUM(( GND ) + ( Xd_0__inst_mult_5_534  ) + ( Xd_0__inst_mult_5_533  ))
// Xd_0__inst_mult_9_545  = CARRY(( GND ) + ( Xd_0__inst_mult_5_534  ) + ( Xd_0__inst_mult_5_533  ))
// Xd_0__inst_mult_9_546  = SHARE(VCC)

	.dataa(!din_a[110]),
	.datab(!din_b[115]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_533 ),
	.sharein(Xd_0__inst_mult_5_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_544 ),
	.cout(Xd_0__inst_mult_9_545 ),
	.shareout(Xd_0__inst_mult_9_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_161 (
// Equation(s):
// Xd_0__inst_mult_2_544  = SUM(( (din_a[32] & din_b[31]) ) + ( Xd_0__inst_mult_2_530  ) + ( Xd_0__inst_mult_2_529  ))
// Xd_0__inst_mult_2_545  = CARRY(( (din_a[32] & din_b[31]) ) + ( Xd_0__inst_mult_2_530  ) + ( Xd_0__inst_mult_2_529  ))
// Xd_0__inst_mult_2_546  = SHARE((din_b[31] & din_a[33]))

	.dataa(!din_a[32]),
	.datab(!din_b[31]),
	.datac(!din_a[33]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_529 ),
	.sharein(Xd_0__inst_mult_2_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_544 ),
	.cout(Xd_0__inst_mult_2_545 ),
	.shareout(Xd_0__inst_mult_2_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_162 (
// Equation(s):
// Xd_0__inst_mult_2_548  = SUM(( (!din_a[31] & (((din_a[30] & din_b[33])))) # (din_a[31] & (!din_b[32] $ (((!din_a[30]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_2_534  ) + ( Xd_0__inst_mult_2_533  ))
// Xd_0__inst_mult_2_549  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[33])))) # (din_a[31] & (!din_b[32] $ (((!din_a[30]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_2_534  ) + ( Xd_0__inst_mult_2_533  ))
// Xd_0__inst_mult_2_550  = SHARE((din_a[31] & (din_b[32] & (din_a[30] & din_b[33]))))

	.dataa(!din_a[31]),
	.datab(!din_b[32]),
	.datac(!din_a[30]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_533 ),
	.sharein(Xd_0__inst_mult_2_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_548 ),
	.cout(Xd_0__inst_mult_2_549 ),
	.shareout(Xd_0__inst_mult_2_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_162 (
// Equation(s):
// Xd_0__inst_mult_13_548  = SUM(( GND ) + ( Xd_0__inst_mult_2_538  ) + ( Xd_0__inst_mult_2_537  ))
// Xd_0__inst_mult_13_549  = CARRY(( GND ) + ( Xd_0__inst_mult_2_538  ) + ( Xd_0__inst_mult_2_537  ))
// Xd_0__inst_mult_13_550  = SHARE(VCC)

	.dataa(!din_a[158]),
	.datab(!din_b[163]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_537 ),
	.sharein(Xd_0__inst_mult_2_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_548 ),
	.cout(Xd_0__inst_mult_13_549 ),
	.shareout(Xd_0__inst_mult_13_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_157 (
// Equation(s):
// Xd_0__inst_mult_3_540  = SUM(( (din_a[44] & din_b[43]) ) + ( Xd_0__inst_mult_3_526  ) + ( Xd_0__inst_mult_3_525  ))
// Xd_0__inst_mult_3_541  = CARRY(( (din_a[44] & din_b[43]) ) + ( Xd_0__inst_mult_3_526  ) + ( Xd_0__inst_mult_3_525  ))
// Xd_0__inst_mult_3_542  = SHARE((din_b[43] & din_a[45]))

	.dataa(!din_a[44]),
	.datab(!din_b[43]),
	.datac(!din_a[45]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_525 ),
	.sharein(Xd_0__inst_mult_3_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_540 ),
	.cout(Xd_0__inst_mult_3_541 ),
	.shareout(Xd_0__inst_mult_3_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_158 (
// Equation(s):
// Xd_0__inst_mult_3_544  = SUM(( (!din_a[43] & (((din_a[42] & din_b[45])))) # (din_a[43] & (!din_b[44] $ (((!din_a[42]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_3_530  ) + ( Xd_0__inst_mult_3_529  ))
// Xd_0__inst_mult_3_545  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[45])))) # (din_a[43] & (!din_b[44] $ (((!din_a[42]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_3_530  ) + ( Xd_0__inst_mult_3_529  ))
// Xd_0__inst_mult_3_546  = SHARE((din_a[43] & (din_b[44] & (din_a[42] & din_b[45]))))

	.dataa(!din_a[43]),
	.datab(!din_b[44]),
	.datac(!din_a[42]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_529 ),
	.sharein(Xd_0__inst_mult_3_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_544 ),
	.cout(Xd_0__inst_mult_3_545 ),
	.shareout(Xd_0__inst_mult_3_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_162 (
// Equation(s):
// Xd_0__inst_mult_8_548  = SUM(( GND ) + ( Xd_0__inst_mult_3_534  ) + ( Xd_0__inst_mult_3_533  ))
// Xd_0__inst_mult_8_549  = CARRY(( GND ) + ( Xd_0__inst_mult_3_534  ) + ( Xd_0__inst_mult_3_533  ))
// Xd_0__inst_mult_8_550  = SHARE(VCC)

	.dataa(!din_a[98]),
	.datab(!din_b[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_533 ),
	.sharein(Xd_0__inst_mult_3_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_548 ),
	.cout(Xd_0__inst_mult_8_549 ),
	.shareout(Xd_0__inst_mult_8_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_161 (
// Equation(s):
// Xd_0__inst_mult_0_544  = SUM(( (din_a[8] & din_b[7]) ) + ( Xd_0__inst_mult_0_530  ) + ( Xd_0__inst_mult_0_529  ))
// Xd_0__inst_mult_0_545  = CARRY(( (din_a[8] & din_b[7]) ) + ( Xd_0__inst_mult_0_530  ) + ( Xd_0__inst_mult_0_529  ))
// Xd_0__inst_mult_0_546  = SHARE((din_b[7] & din_a[9]))

	.dataa(!din_a[8]),
	.datab(!din_b[7]),
	.datac(!din_a[9]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_529 ),
	.sharein(Xd_0__inst_mult_0_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_544 ),
	.cout(Xd_0__inst_mult_0_545 ),
	.shareout(Xd_0__inst_mult_0_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_162 (
// Equation(s):
// Xd_0__inst_mult_0_548  = SUM(( (!din_a[7] & (((din_a[6] & din_b[9])))) # (din_a[7] & (!din_b[8] $ (((!din_a[6]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_0_534  ) + ( Xd_0__inst_mult_0_533  ))
// Xd_0__inst_mult_0_549  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[9])))) # (din_a[7] & (!din_b[8] $ (((!din_a[6]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_0_534  ) + ( Xd_0__inst_mult_0_533  ))
// Xd_0__inst_mult_0_550  = SHARE((din_a[7] & (din_b[8] & (din_a[6] & din_b[9]))))

	.dataa(!din_a[7]),
	.datab(!din_b[8]),
	.datac(!din_a[6]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_533 ),
	.sharein(Xd_0__inst_mult_0_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_548 ),
	.cout(Xd_0__inst_mult_0_549 ),
	.shareout(Xd_0__inst_mult_0_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_162 (
// Equation(s):
// Xd_0__inst_mult_11_548  = SUM(( GND ) + ( Xd_0__inst_mult_0_538  ) + ( Xd_0__inst_mult_0_537  ))
// Xd_0__inst_mult_11_549  = CARRY(( GND ) + ( Xd_0__inst_mult_0_538  ) + ( Xd_0__inst_mult_0_537  ))
// Xd_0__inst_mult_11_550  = SHARE(VCC)

	.dataa(!din_a[134]),
	.datab(!din_b[139]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_537 ),
	.sharein(Xd_0__inst_mult_0_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_548 ),
	.cout(Xd_0__inst_mult_11_549 ),
	.shareout(Xd_0__inst_mult_11_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_162 (
// Equation(s):
// Xd_0__inst_mult_1_548  = SUM(( (din_a[20] & din_b[19]) ) + ( Xd_0__inst_mult_1_530  ) + ( Xd_0__inst_mult_1_529  ))
// Xd_0__inst_mult_1_549  = CARRY(( (din_a[20] & din_b[19]) ) + ( Xd_0__inst_mult_1_530  ) + ( Xd_0__inst_mult_1_529  ))
// Xd_0__inst_mult_1_550  = SHARE((din_b[19] & din_a[21]))

	.dataa(!din_a[20]),
	.datab(!din_b[19]),
	.datac(!din_a[21]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_529 ),
	.sharein(Xd_0__inst_mult_1_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_548 ),
	.cout(Xd_0__inst_mult_1_549 ),
	.shareout(Xd_0__inst_mult_1_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_163 (
// Equation(s):
// Xd_0__inst_mult_1_552  = SUM(( (!din_a[19] & (((din_a[18] & din_b[21])))) # (din_a[19] & (!din_b[20] $ (((!din_a[18]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_1_534  ) + ( Xd_0__inst_mult_1_533  ))
// Xd_0__inst_mult_1_553  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[21])))) # (din_a[19] & (!din_b[20] $ (((!din_a[18]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_1_534  ) + ( Xd_0__inst_mult_1_533  ))
// Xd_0__inst_mult_1_554  = SHARE((din_a[19] & (din_b[20] & (din_a[18] & din_b[21]))))

	.dataa(!din_a[19]),
	.datab(!din_b[20]),
	.datac(!din_a[18]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_533 ),
	.sharein(Xd_0__inst_mult_1_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_552 ),
	.cout(Xd_0__inst_mult_1_553 ),
	.shareout(Xd_0__inst_mult_1_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_158 (
// Equation(s):
// Xd_0__inst_mult_10_544  = SUM(( GND ) + ( Xd_0__inst_mult_1_538  ) + ( Xd_0__inst_mult_1_537  ))
// Xd_0__inst_mult_10_545  = CARRY(( GND ) + ( Xd_0__inst_mult_1_538  ) + ( Xd_0__inst_mult_1_537  ))
// Xd_0__inst_mult_10_546  = SHARE(VCC)

	.dataa(!din_a[122]),
	.datab(!din_b[127]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_537 ),
	.sharein(Xd_0__inst_mult_1_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_544 ),
	.cout(Xd_0__inst_mult_10_545 ),
	.shareout(Xd_0__inst_mult_10_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_162 (
// Equation(s):
// Xd_0__inst_mult_12_560  = SUM(( (din_a[152] & din_b[152]) ) + ( Xd_0__inst_mult_12_558  ) + ( Xd_0__inst_mult_12_557  ))
// Xd_0__inst_mult_12_561  = CARRY(( (din_a[152] & din_b[152]) ) + ( Xd_0__inst_mult_12_558  ) + ( Xd_0__inst_mult_12_557  ))
// Xd_0__inst_mult_12_562  = SHARE(GND)

	.dataa(!din_a[152]),
	.datab(!din_b[152]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_557 ),
	.sharein(Xd_0__inst_mult_12_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_560 ),
	.cout(Xd_0__inst_mult_12_561 ),
	.shareout(Xd_0__inst_mult_12_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_163 (
// Equation(s):
// Xd_0__inst_mult_13_552  = SUM(( (din_a[164] & din_b[164]) ) + ( Xd_0__inst_mult_13_542  ) + ( Xd_0__inst_mult_13_541  ))
// Xd_0__inst_mult_13_553  = CARRY(( (din_a[164] & din_b[164]) ) + ( Xd_0__inst_mult_13_542  ) + ( Xd_0__inst_mult_13_541  ))
// Xd_0__inst_mult_13_554  = SHARE(GND)

	.dataa(!din_a[164]),
	.datab(!din_b[164]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_541 ),
	.sharein(Xd_0__inst_mult_13_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_552 ),
	.cout(Xd_0__inst_mult_13_553 ),
	.shareout(Xd_0__inst_mult_13_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_164 (
// Equation(s):
// Xd_0__inst_mult_13_556  = SUM(( (!din_a[163] & (((din_a[162] & din_b[166])))) # (din_a[163] & (!din_b[165] $ (((!din_a[162]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_13_546  ) + ( Xd_0__inst_mult_13_545  ))
// Xd_0__inst_mult_13_557  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[166])))) # (din_a[163] & (!din_b[165] $ (((!din_a[162]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_13_546  ) + ( Xd_0__inst_mult_13_545  ))
// Xd_0__inst_mult_13_558  = SHARE((din_a[163] & (din_b[165] & (din_a[162] & din_b[166]))))

	.dataa(!din_a[163]),
	.datab(!din_b[165]),
	.datac(!din_a[162]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_545 ),
	.sharein(Xd_0__inst_mult_13_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_556 ),
	.cout(Xd_0__inst_mult_13_557 ),
	.shareout(Xd_0__inst_mult_13_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_164 (
// Equation(s):
// Xd_0__inst_mult_14_556  = SUM(( (din_a[176] & din_b[176]) ) + ( Xd_0__inst_mult_14_546  ) + ( Xd_0__inst_mult_14_545  ))
// Xd_0__inst_mult_14_557  = CARRY(( (din_a[176] & din_b[176]) ) + ( Xd_0__inst_mult_14_546  ) + ( Xd_0__inst_mult_14_545  ))
// Xd_0__inst_mult_14_558  = SHARE(GND)

	.dataa(!din_a[176]),
	.datab(!din_b[176]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_545 ),
	.sharein(Xd_0__inst_mult_14_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_556 ),
	.cout(Xd_0__inst_mult_14_557 ),
	.shareout(Xd_0__inst_mult_14_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_165 (
// Equation(s):
// Xd_0__inst_mult_14_560  = SUM(( (!din_a[175] & (((din_a[174] & din_b[178])))) # (din_a[175] & (!din_b[177] $ (((!din_a[174]) # (!din_b[178]))))) ) + ( Xd_0__inst_mult_14_550  ) + ( Xd_0__inst_mult_14_549  ))
// Xd_0__inst_mult_14_561  = CARRY(( (!din_a[175] & (((din_a[174] & din_b[178])))) # (din_a[175] & (!din_b[177] $ (((!din_a[174]) # (!din_b[178]))))) ) + ( Xd_0__inst_mult_14_550  ) + ( Xd_0__inst_mult_14_549  ))
// Xd_0__inst_mult_14_562  = SHARE((din_a[175] & (din_b[177] & (din_a[174] & din_b[178]))))

	.dataa(!din_a[175]),
	.datab(!din_b[177]),
	.datac(!din_a[174]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_549 ),
	.sharein(Xd_0__inst_mult_14_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_560 ),
	.cout(Xd_0__inst_mult_14_561 ),
	.shareout(Xd_0__inst_mult_14_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_167 (
// Equation(s):
// Xd_0__inst_mult_15_568  = SUM(( (din_a[188] & din_b[188]) ) + ( Xd_0__inst_mult_15_566  ) + ( Xd_0__inst_mult_15_565  ))
// Xd_0__inst_mult_15_569  = CARRY(( (din_a[188] & din_b[188]) ) + ( Xd_0__inst_mult_15_566  ) + ( Xd_0__inst_mult_15_565  ))
// Xd_0__inst_mult_15_570  = SHARE(GND)

	.dataa(!din_a[188]),
	.datab(!din_b[188]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_565 ),
	.sharein(Xd_0__inst_mult_15_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_568 ),
	.cout(Xd_0__inst_mult_15_569 ),
	.shareout(Xd_0__inst_mult_15_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_159 (
// Equation(s):
// Xd_0__inst_mult_10_548  = SUM(( (din_a[128] & din_b[128]) ) + ( Xd_0__inst_mult_10_538  ) + ( Xd_0__inst_mult_10_537  ))
// Xd_0__inst_mult_10_549  = CARRY(( (din_a[128] & din_b[128]) ) + ( Xd_0__inst_mult_10_538  ) + ( Xd_0__inst_mult_10_537  ))
// Xd_0__inst_mult_10_550  = SHARE(GND)

	.dataa(!din_a[128]),
	.datab(!din_b[128]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_537 ),
	.sharein(Xd_0__inst_mult_10_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_548 ),
	.cout(Xd_0__inst_mult_10_549 ),
	.shareout(Xd_0__inst_mult_10_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_160 (
// Equation(s):
// Xd_0__inst_mult_10_552  = SUM(( (!din_a[127] & (((din_a[126] & din_b[130])))) # (din_a[127] & (!din_b[129] $ (((!din_a[126]) # (!din_b[130]))))) ) + ( Xd_0__inst_mult_10_542  ) + ( Xd_0__inst_mult_10_541  ))
// Xd_0__inst_mult_10_553  = CARRY(( (!din_a[127] & (((din_a[126] & din_b[130])))) # (din_a[127] & (!din_b[129] $ (((!din_a[126]) # (!din_b[130]))))) ) + ( Xd_0__inst_mult_10_542  ) + ( Xd_0__inst_mult_10_541  ))
// Xd_0__inst_mult_10_554  = SHARE((din_a[127] & (din_b[129] & (din_a[126] & din_b[130]))))

	.dataa(!din_a[127]),
	.datab(!din_b[129]),
	.datac(!din_a[126]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_541 ),
	.sharein(Xd_0__inst_mult_10_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_552 ),
	.cout(Xd_0__inst_mult_10_553 ),
	.shareout(Xd_0__inst_mult_10_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_163 (
// Equation(s):
// Xd_0__inst_mult_11_552  = SUM(( (din_a[140] & din_b[140]) ) + ( Xd_0__inst_mult_11_542  ) + ( Xd_0__inst_mult_11_541  ))
// Xd_0__inst_mult_11_553  = CARRY(( (din_a[140] & din_b[140]) ) + ( Xd_0__inst_mult_11_542  ) + ( Xd_0__inst_mult_11_541  ))
// Xd_0__inst_mult_11_554  = SHARE(GND)

	.dataa(!din_a[140]),
	.datab(!din_b[140]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_541 ),
	.sharein(Xd_0__inst_mult_11_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_552 ),
	.cout(Xd_0__inst_mult_11_553 ),
	.shareout(Xd_0__inst_mult_11_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_164 (
// Equation(s):
// Xd_0__inst_mult_11_556  = SUM(( (!din_a[139] & (((din_a[138] & din_b[142])))) # (din_a[139] & (!din_b[141] $ (((!din_a[138]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_11_546  ) + ( Xd_0__inst_mult_11_545  ))
// Xd_0__inst_mult_11_557  = CARRY(( (!din_a[139] & (((din_a[138] & din_b[142])))) # (din_a[139] & (!din_b[141] $ (((!din_a[138]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_11_546  ) + ( Xd_0__inst_mult_11_545  ))
// Xd_0__inst_mult_11_558  = SHARE((din_a[139] & (din_b[141] & (din_a[138] & din_b[142]))))

	.dataa(!din_a[139]),
	.datab(!din_b[141]),
	.datac(!din_a[138]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_545 ),
	.sharein(Xd_0__inst_mult_11_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_556 ),
	.cout(Xd_0__inst_mult_11_557 ),
	.shareout(Xd_0__inst_mult_11_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_163 (
// Equation(s):
// Xd_0__inst_mult_8_552  = SUM(( (din_a[104] & din_b[104]) ) + ( Xd_0__inst_mult_8_542  ) + ( Xd_0__inst_mult_8_541  ))
// Xd_0__inst_mult_8_553  = CARRY(( (din_a[104] & din_b[104]) ) + ( Xd_0__inst_mult_8_542  ) + ( Xd_0__inst_mult_8_541  ))
// Xd_0__inst_mult_8_554  = SHARE(GND)

	.dataa(!din_a[104]),
	.datab(!din_b[104]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_541 ),
	.sharein(Xd_0__inst_mult_8_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_552 ),
	.cout(Xd_0__inst_mult_8_553 ),
	.shareout(Xd_0__inst_mult_8_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_164 (
// Equation(s):
// Xd_0__inst_mult_8_556  = SUM(( (!din_a[103] & (((din_a[102] & din_b[106])))) # (din_a[103] & (!din_b[105] $ (((!din_a[102]) # (!din_b[106]))))) ) + ( Xd_0__inst_mult_8_546  ) + ( Xd_0__inst_mult_8_545  ))
// Xd_0__inst_mult_8_557  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[106])))) # (din_a[103] & (!din_b[105] $ (((!din_a[102]) # (!din_b[106]))))) ) + ( Xd_0__inst_mult_8_546  ) + ( Xd_0__inst_mult_8_545  ))
// Xd_0__inst_mult_8_558  = SHARE((din_a[103] & (din_b[105] & (din_a[102] & din_b[106]))))

	.dataa(!din_a[103]),
	.datab(!din_b[105]),
	.datac(!din_a[102]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_545 ),
	.sharein(Xd_0__inst_mult_8_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_556 ),
	.cout(Xd_0__inst_mult_8_557 ),
	.shareout(Xd_0__inst_mult_8_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_159 (
// Equation(s):
// Xd_0__inst_mult_9_548  = SUM(( (din_a[116] & din_b[116]) ) + ( Xd_0__inst_mult_9_538  ) + ( Xd_0__inst_mult_9_537  ))
// Xd_0__inst_mult_9_549  = CARRY(( (din_a[116] & din_b[116]) ) + ( Xd_0__inst_mult_9_538  ) + ( Xd_0__inst_mult_9_537  ))
// Xd_0__inst_mult_9_550  = SHARE(GND)

	.dataa(!din_a[116]),
	.datab(!din_b[116]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_537 ),
	.sharein(Xd_0__inst_mult_9_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_548 ),
	.cout(Xd_0__inst_mult_9_549 ),
	.shareout(Xd_0__inst_mult_9_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_160 (
// Equation(s):
// Xd_0__inst_mult_9_552  = SUM(( (!din_a[115] & (((din_a[114] & din_b[118])))) # (din_a[115] & (!din_b[117] $ (((!din_a[114]) # (!din_b[118]))))) ) + ( Xd_0__inst_mult_9_542  ) + ( Xd_0__inst_mult_9_541  ))
// Xd_0__inst_mult_9_553  = CARRY(( (!din_a[115] & (((din_a[114] & din_b[118])))) # (din_a[115] & (!din_b[117] $ (((!din_a[114]) # (!din_b[118]))))) ) + ( Xd_0__inst_mult_9_542  ) + ( Xd_0__inst_mult_9_541  ))
// Xd_0__inst_mult_9_554  = SHARE((din_a[115] & (din_b[117] & (din_a[114] & din_b[118]))))

	.dataa(!din_a[115]),
	.datab(!din_b[117]),
	.datac(!din_a[114]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_541 ),
	.sharein(Xd_0__inst_mult_9_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_552 ),
	.cout(Xd_0__inst_mult_9_553 ),
	.shareout(Xd_0__inst_mult_9_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_159 (
// Equation(s):
// Xd_0__inst_mult_6_548  = SUM(( (din_a[80] & din_b[80]) ) + ( Xd_0__inst_mult_6_538  ) + ( Xd_0__inst_mult_6_537  ))
// Xd_0__inst_mult_6_549  = CARRY(( (din_a[80] & din_b[80]) ) + ( Xd_0__inst_mult_6_538  ) + ( Xd_0__inst_mult_6_537  ))
// Xd_0__inst_mult_6_550  = SHARE(GND)

	.dataa(!din_a[80]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_537 ),
	.sharein(Xd_0__inst_mult_6_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_548 ),
	.cout(Xd_0__inst_mult_6_549 ),
	.shareout(Xd_0__inst_mult_6_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_160 (
// Equation(s):
// Xd_0__inst_mult_6_552  = SUM(( (!din_a[79] & (((din_a[78] & din_b[82])))) # (din_a[79] & (!din_b[81] $ (((!din_a[78]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_542  ) + ( Xd_0__inst_mult_6_541  ))
// Xd_0__inst_mult_6_553  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[82])))) # (din_a[79] & (!din_b[81] $ (((!din_a[78]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_542  ) + ( Xd_0__inst_mult_6_541  ))
// Xd_0__inst_mult_6_554  = SHARE((din_a[79] & (din_b[81] & (din_a[78] & din_b[82]))))

	.dataa(!din_a[79]),
	.datab(!din_b[81]),
	.datac(!din_a[78]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_541 ),
	.sharein(Xd_0__inst_mult_6_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_552 ),
	.cout(Xd_0__inst_mult_6_553 ),
	.shareout(Xd_0__inst_mult_6_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_159 (
// Equation(s):
// Xd_0__inst_mult_7_548  = SUM(( (din_a[92] & din_b[92]) ) + ( Xd_0__inst_mult_7_538  ) + ( Xd_0__inst_mult_7_537  ))
// Xd_0__inst_mult_7_549  = CARRY(( (din_a[92] & din_b[92]) ) + ( Xd_0__inst_mult_7_538  ) + ( Xd_0__inst_mult_7_537  ))
// Xd_0__inst_mult_7_550  = SHARE(GND)

	.dataa(!din_a[92]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_537 ),
	.sharein(Xd_0__inst_mult_7_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_548 ),
	.cout(Xd_0__inst_mult_7_549 ),
	.shareout(Xd_0__inst_mult_7_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_160 (
// Equation(s):
// Xd_0__inst_mult_7_552  = SUM(( (!din_a[91] & (((din_a[90] & din_b[94])))) # (din_a[91] & (!din_b[93] $ (((!din_a[90]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_542  ) + ( Xd_0__inst_mult_7_541  ))
// Xd_0__inst_mult_7_553  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[94])))) # (din_a[91] & (!din_b[93] $ (((!din_a[90]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_542  ) + ( Xd_0__inst_mult_7_541  ))
// Xd_0__inst_mult_7_554  = SHARE((din_a[91] & (din_b[93] & (din_a[90] & din_b[94]))))

	.dataa(!din_a[91]),
	.datab(!din_b[93]),
	.datac(!din_a[90]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_541 ),
	.sharein(Xd_0__inst_mult_7_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_552 ),
	.cout(Xd_0__inst_mult_7_553 ),
	.shareout(Xd_0__inst_mult_7_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_166 (
// Equation(s):
// Xd_0__inst_mult_4_564  = SUM(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_4_562  ) + ( Xd_0__inst_mult_4_561  ))
// Xd_0__inst_mult_4_565  = CARRY(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_4_562  ) + ( Xd_0__inst_mult_4_561  ))
// Xd_0__inst_mult_4_566  = SHARE(GND)

	.dataa(!din_a[56]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_561 ),
	.sharein(Xd_0__inst_mult_4_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_564 ),
	.cout(Xd_0__inst_mult_4_565 ),
	.shareout(Xd_0__inst_mult_4_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_159 (
// Equation(s):
// Xd_0__inst_mult_5_548  = SUM(( (din_a[68] & din_b[68]) ) + ( Xd_0__inst_mult_5_542  ) + ( Xd_0__inst_mult_5_541  ))
// Xd_0__inst_mult_5_549  = CARRY(( (din_a[68] & din_b[68]) ) + ( Xd_0__inst_mult_5_542  ) + ( Xd_0__inst_mult_5_541  ))
// Xd_0__inst_mult_5_550  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_541 ),
	.sharein(Xd_0__inst_mult_5_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_548 ),
	.cout(Xd_0__inst_mult_5_549 ),
	.shareout(Xd_0__inst_mult_5_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_160 (
// Equation(s):
// Xd_0__inst_mult_5_552  = SUM(( (!din_a[67] & (((din_a[66] & din_b[70])))) # (din_a[67] & (!din_b[69] $ (((!din_a[66]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_546  ) + ( Xd_0__inst_mult_5_545  ))
// Xd_0__inst_mult_5_553  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[70])))) # (din_a[67] & (!din_b[69] $ (((!din_a[66]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_546  ) + ( Xd_0__inst_mult_5_545  ))
// Xd_0__inst_mult_5_554  = SHARE((din_a[67] & (din_b[69] & (din_a[66] & din_b[70]))))

	.dataa(!din_a[67]),
	.datab(!din_b[69]),
	.datac(!din_a[66]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_545 ),
	.sharein(Xd_0__inst_mult_5_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_552 ),
	.cout(Xd_0__inst_mult_5_553 ),
	.shareout(Xd_0__inst_mult_5_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_163 (
// Equation(s):
// Xd_0__inst_mult_2_552  = SUM(( (din_a[32] & din_b[32]) ) + ( Xd_0__inst_mult_2_546  ) + ( Xd_0__inst_mult_2_545  ))
// Xd_0__inst_mult_2_553  = CARRY(( (din_a[32] & din_b[32]) ) + ( Xd_0__inst_mult_2_546  ) + ( Xd_0__inst_mult_2_545  ))
// Xd_0__inst_mult_2_554  = SHARE(GND)

	.dataa(!din_a[32]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_545 ),
	.sharein(Xd_0__inst_mult_2_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_552 ),
	.cout(Xd_0__inst_mult_2_553 ),
	.shareout(Xd_0__inst_mult_2_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_164 (
// Equation(s):
// Xd_0__inst_mult_2_556  = SUM(( (!din_a[31] & (((din_a[30] & din_b[34])))) # (din_a[31] & (!din_b[33] $ (((!din_a[30]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_550  ) + ( Xd_0__inst_mult_2_549  ))
// Xd_0__inst_mult_2_557  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[34])))) # (din_a[31] & (!din_b[33] $ (((!din_a[30]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_550  ) + ( Xd_0__inst_mult_2_549  ))
// Xd_0__inst_mult_2_558  = SHARE((din_a[31] & (din_b[33] & (din_a[30] & din_b[34]))))

	.dataa(!din_a[31]),
	.datab(!din_b[33]),
	.datac(!din_a[30]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_549 ),
	.sharein(Xd_0__inst_mult_2_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_556 ),
	.cout(Xd_0__inst_mult_2_557 ),
	.shareout(Xd_0__inst_mult_2_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_159 (
// Equation(s):
// Xd_0__inst_mult_3_548  = SUM(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_3_542  ) + ( Xd_0__inst_mult_3_541  ))
// Xd_0__inst_mult_3_549  = CARRY(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_3_542  ) + ( Xd_0__inst_mult_3_541  ))
// Xd_0__inst_mult_3_550  = SHARE(GND)

	.dataa(!din_a[44]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_541 ),
	.sharein(Xd_0__inst_mult_3_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_548 ),
	.cout(Xd_0__inst_mult_3_549 ),
	.shareout(Xd_0__inst_mult_3_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_160 (
// Equation(s):
// Xd_0__inst_mult_3_552  = SUM(( (!din_a[43] & (((din_a[42] & din_b[46])))) # (din_a[43] & (!din_b[45] $ (((!din_a[42]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_546  ) + ( Xd_0__inst_mult_3_545  ))
// Xd_0__inst_mult_3_553  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[46])))) # (din_a[43] & (!din_b[45] $ (((!din_a[42]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_546  ) + ( Xd_0__inst_mult_3_545  ))
// Xd_0__inst_mult_3_554  = SHARE((din_a[43] & (din_b[45] & (din_a[42] & din_b[46]))))

	.dataa(!din_a[43]),
	.datab(!din_b[45]),
	.datac(!din_a[42]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_545 ),
	.sharein(Xd_0__inst_mult_3_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_552 ),
	.cout(Xd_0__inst_mult_3_553 ),
	.shareout(Xd_0__inst_mult_3_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_163 (
// Equation(s):
// Xd_0__inst_mult_0_552  = SUM(( (din_a[8] & din_b[8]) ) + ( Xd_0__inst_mult_0_546  ) + ( Xd_0__inst_mult_0_545  ))
// Xd_0__inst_mult_0_553  = CARRY(( (din_a[8] & din_b[8]) ) + ( Xd_0__inst_mult_0_546  ) + ( Xd_0__inst_mult_0_545  ))
// Xd_0__inst_mult_0_554  = SHARE(GND)

	.dataa(!din_a[8]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_545 ),
	.sharein(Xd_0__inst_mult_0_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_552 ),
	.cout(Xd_0__inst_mult_0_553 ),
	.shareout(Xd_0__inst_mult_0_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_164 (
// Equation(s):
// Xd_0__inst_mult_0_556  = SUM(( (!din_a[7] & (((din_a[6] & din_b[10])))) # (din_a[7] & (!din_b[9] $ (((!din_a[6]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_550  ) + ( Xd_0__inst_mult_0_549  ))
// Xd_0__inst_mult_0_557  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[10])))) # (din_a[7] & (!din_b[9] $ (((!din_a[6]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_550  ) + ( Xd_0__inst_mult_0_549  ))
// Xd_0__inst_mult_0_558  = SHARE((din_a[7] & (din_b[9] & (din_a[6] & din_b[10]))))

	.dataa(!din_a[7]),
	.datab(!din_b[9]),
	.datac(!din_a[6]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_549 ),
	.sharein(Xd_0__inst_mult_0_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_556 ),
	.cout(Xd_0__inst_mult_0_557 ),
	.shareout(Xd_0__inst_mult_0_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_164 (
// Equation(s):
// Xd_0__inst_mult_1_556  = SUM(( (din_a[20] & din_b[20]) ) + ( Xd_0__inst_mult_1_550  ) + ( Xd_0__inst_mult_1_549  ))
// Xd_0__inst_mult_1_557  = CARRY(( (din_a[20] & din_b[20]) ) + ( Xd_0__inst_mult_1_550  ) + ( Xd_0__inst_mult_1_549  ))
// Xd_0__inst_mult_1_558  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_549 ),
	.sharein(Xd_0__inst_mult_1_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_556 ),
	.cout(Xd_0__inst_mult_1_557 ),
	.shareout(Xd_0__inst_mult_1_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_165 (
// Equation(s):
// Xd_0__inst_mult_1_560  = SUM(( (!din_a[19] & (((din_a[18] & din_b[22])))) # (din_a[19] & (!din_b[21] $ (((!din_a[18]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_554  ) + ( Xd_0__inst_mult_1_553  ))
// Xd_0__inst_mult_1_561  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[22])))) # (din_a[19] & (!din_b[21] $ (((!din_a[18]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_554  ) + ( Xd_0__inst_mult_1_553  ))
// Xd_0__inst_mult_1_562  = SHARE((din_a[19] & (din_b[21] & (din_a[18] & din_b[22]))))

	.dataa(!din_a[19]),
	.datab(!din_b[21]),
	.datac(!din_a[18]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_553 ),
	.sharein(Xd_0__inst_mult_1_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_560 ),
	.cout(Xd_0__inst_mult_1_561 ),
	.shareout(Xd_0__inst_mult_1_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_163 (
// Equation(s):
// Xd_0__inst_mult_12_564  = SUM(( GND ) + ( Xd_0__inst_mult_12_562  ) + ( Xd_0__inst_mult_12_561  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_561 ),
	.sharein(Xd_0__inst_mult_12_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_564 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_165 (
// Equation(s):
// Xd_0__inst_mult_13_560  = SUM(( GND ) + ( Xd_0__inst_mult_13_554  ) + ( Xd_0__inst_mult_13_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_553 ),
	.sharein(Xd_0__inst_mult_13_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_166 (
// Equation(s):
// Xd_0__inst_mult_13_564  = SUM(( (!din_a[164] & (((din_a[163] & din_b[166])))) # (din_a[164] & (!din_b[165] $ (((!din_a[163]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_13_558  ) + ( Xd_0__inst_mult_13_557  ))
// Xd_0__inst_mult_13_565  = CARRY(( (!din_a[164] & (((din_a[163] & din_b[166])))) # (din_a[164] & (!din_b[165] $ (((!din_a[163]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_13_558  ) + ( Xd_0__inst_mult_13_557  ))
// Xd_0__inst_mult_13_566  = SHARE((din_a[164] & (din_b[165] & (din_a[163] & din_b[166]))))

	.dataa(!din_a[164]),
	.datab(!din_b[165]),
	.datac(!din_a[163]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_557 ),
	.sharein(Xd_0__inst_mult_13_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_564 ),
	.cout(Xd_0__inst_mult_13_565 ),
	.shareout(Xd_0__inst_mult_13_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_166 (
// Equation(s):
// Xd_0__inst_mult_14_564  = SUM(( GND ) + ( Xd_0__inst_mult_14_558  ) + ( Xd_0__inst_mult_14_557  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_557 ),
	.sharein(Xd_0__inst_mult_14_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_564 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_167 (
// Equation(s):
// Xd_0__inst_mult_14_568  = SUM(( (!din_a[176] & (((din_a[175] & din_b[178])))) # (din_a[176] & (!din_b[177] $ (((!din_a[175]) # (!din_b[178]))))) ) + ( Xd_0__inst_mult_14_562  ) + ( Xd_0__inst_mult_14_561  ))
// Xd_0__inst_mult_14_569  = CARRY(( (!din_a[176] & (((din_a[175] & din_b[178])))) # (din_a[176] & (!din_b[177] $ (((!din_a[175]) # (!din_b[178]))))) ) + ( Xd_0__inst_mult_14_562  ) + ( Xd_0__inst_mult_14_561  ))
// Xd_0__inst_mult_14_570  = SHARE((din_a[176] & (din_b[177] & (din_a[175] & din_b[178]))))

	.dataa(!din_a[176]),
	.datab(!din_b[177]),
	.datac(!din_a[175]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_561 ),
	.sharein(Xd_0__inst_mult_14_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_568 ),
	.cout(Xd_0__inst_mult_14_569 ),
	.shareout(Xd_0__inst_mult_14_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_168 (
// Equation(s):
// Xd_0__inst_mult_15_572  = SUM(( GND ) + ( Xd_0__inst_mult_15_570  ) + ( Xd_0__inst_mult_15_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_569 ),
	.sharein(Xd_0__inst_mult_15_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_161 (
// Equation(s):
// Xd_0__inst_mult_10_556  = SUM(( GND ) + ( Xd_0__inst_mult_10_550  ) + ( Xd_0__inst_mult_10_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_549 ),
	.sharein(Xd_0__inst_mult_10_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_162 (
// Equation(s):
// Xd_0__inst_mult_10_560  = SUM(( (!din_a[128] & (((din_a[127] & din_b[130])))) # (din_a[128] & (!din_b[129] $ (((!din_a[127]) # (!din_b[130]))))) ) + ( Xd_0__inst_mult_10_554  ) + ( Xd_0__inst_mult_10_553  ))
// Xd_0__inst_mult_10_561  = CARRY(( (!din_a[128] & (((din_a[127] & din_b[130])))) # (din_a[128] & (!din_b[129] $ (((!din_a[127]) # (!din_b[130]))))) ) + ( Xd_0__inst_mult_10_554  ) + ( Xd_0__inst_mult_10_553  ))
// Xd_0__inst_mult_10_562  = SHARE((din_a[128] & (din_b[129] & (din_a[127] & din_b[130]))))

	.dataa(!din_a[128]),
	.datab(!din_b[129]),
	.datac(!din_a[127]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_553 ),
	.sharein(Xd_0__inst_mult_10_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_560 ),
	.cout(Xd_0__inst_mult_10_561 ),
	.shareout(Xd_0__inst_mult_10_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_165 (
// Equation(s):
// Xd_0__inst_mult_11_560  = SUM(( GND ) + ( Xd_0__inst_mult_11_554  ) + ( Xd_0__inst_mult_11_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_553 ),
	.sharein(Xd_0__inst_mult_11_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_166 (
// Equation(s):
// Xd_0__inst_mult_11_564  = SUM(( (!din_a[140] & (((din_a[139] & din_b[142])))) # (din_a[140] & (!din_b[141] $ (((!din_a[139]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_11_558  ) + ( Xd_0__inst_mult_11_557  ))
// Xd_0__inst_mult_11_565  = CARRY(( (!din_a[140] & (((din_a[139] & din_b[142])))) # (din_a[140] & (!din_b[141] $ (((!din_a[139]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_11_558  ) + ( Xd_0__inst_mult_11_557  ))
// Xd_0__inst_mult_11_566  = SHARE((din_a[140] & (din_b[141] & (din_a[139] & din_b[142]))))

	.dataa(!din_a[140]),
	.datab(!din_b[141]),
	.datac(!din_a[139]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_557 ),
	.sharein(Xd_0__inst_mult_11_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_564 ),
	.cout(Xd_0__inst_mult_11_565 ),
	.shareout(Xd_0__inst_mult_11_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_165 (
// Equation(s):
// Xd_0__inst_mult_8_560  = SUM(( GND ) + ( Xd_0__inst_mult_8_554  ) + ( Xd_0__inst_mult_8_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_553 ),
	.sharein(Xd_0__inst_mult_8_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_166 (
// Equation(s):
// Xd_0__inst_mult_8_564  = SUM(( (!din_a[104] & (((din_a[103] & din_b[106])))) # (din_a[104] & (!din_b[105] $ (((!din_a[103]) # (!din_b[106]))))) ) + ( Xd_0__inst_mult_8_558  ) + ( Xd_0__inst_mult_8_557  ))
// Xd_0__inst_mult_8_565  = CARRY(( (!din_a[104] & (((din_a[103] & din_b[106])))) # (din_a[104] & (!din_b[105] $ (((!din_a[103]) # (!din_b[106]))))) ) + ( Xd_0__inst_mult_8_558  ) + ( Xd_0__inst_mult_8_557  ))
// Xd_0__inst_mult_8_566  = SHARE((din_a[104] & (din_b[105] & (din_a[103] & din_b[106]))))

	.dataa(!din_a[104]),
	.datab(!din_b[105]),
	.datac(!din_a[103]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_557 ),
	.sharein(Xd_0__inst_mult_8_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_564 ),
	.cout(Xd_0__inst_mult_8_565 ),
	.shareout(Xd_0__inst_mult_8_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_161 (
// Equation(s):
// Xd_0__inst_mult_9_556  = SUM(( GND ) + ( Xd_0__inst_mult_9_550  ) + ( Xd_0__inst_mult_9_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_549 ),
	.sharein(Xd_0__inst_mult_9_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_162 (
// Equation(s):
// Xd_0__inst_mult_9_560  = SUM(( (!din_a[116] & (((din_a[115] & din_b[118])))) # (din_a[116] & (!din_b[117] $ (((!din_a[115]) # (!din_b[118]))))) ) + ( Xd_0__inst_mult_9_554  ) + ( Xd_0__inst_mult_9_553  ))
// Xd_0__inst_mult_9_561  = CARRY(( (!din_a[116] & (((din_a[115] & din_b[118])))) # (din_a[116] & (!din_b[117] $ (((!din_a[115]) # (!din_b[118]))))) ) + ( Xd_0__inst_mult_9_554  ) + ( Xd_0__inst_mult_9_553  ))
// Xd_0__inst_mult_9_562  = SHARE((din_a[116] & (din_b[117] & (din_a[115] & din_b[118]))))

	.dataa(!din_a[116]),
	.datab(!din_b[117]),
	.datac(!din_a[115]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_553 ),
	.sharein(Xd_0__inst_mult_9_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_560 ),
	.cout(Xd_0__inst_mult_9_561 ),
	.shareout(Xd_0__inst_mult_9_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_161 (
// Equation(s):
// Xd_0__inst_mult_6_556  = SUM(( GND ) + ( Xd_0__inst_mult_6_550  ) + ( Xd_0__inst_mult_6_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_549 ),
	.sharein(Xd_0__inst_mult_6_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_162 (
// Equation(s):
// Xd_0__inst_mult_6_560  = SUM(( (!din_a[80] & (((din_a[79] & din_b[82])))) # (din_a[80] & (!din_b[81] $ (((!din_a[79]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_554  ) + ( Xd_0__inst_mult_6_553  ))
// Xd_0__inst_mult_6_561  = CARRY(( (!din_a[80] & (((din_a[79] & din_b[82])))) # (din_a[80] & (!din_b[81] $ (((!din_a[79]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_554  ) + ( Xd_0__inst_mult_6_553  ))
// Xd_0__inst_mult_6_562  = SHARE((din_a[80] & (din_b[81] & (din_a[79] & din_b[82]))))

	.dataa(!din_a[80]),
	.datab(!din_b[81]),
	.datac(!din_a[79]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_553 ),
	.sharein(Xd_0__inst_mult_6_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_560 ),
	.cout(Xd_0__inst_mult_6_561 ),
	.shareout(Xd_0__inst_mult_6_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_161 (
// Equation(s):
// Xd_0__inst_mult_7_556  = SUM(( GND ) + ( Xd_0__inst_mult_7_550  ) + ( Xd_0__inst_mult_7_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_549 ),
	.sharein(Xd_0__inst_mult_7_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_162 (
// Equation(s):
// Xd_0__inst_mult_7_560  = SUM(( (!din_a[92] & (((din_a[91] & din_b[94])))) # (din_a[92] & (!din_b[93] $ (((!din_a[91]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_554  ) + ( Xd_0__inst_mult_7_553  ))
// Xd_0__inst_mult_7_561  = CARRY(( (!din_a[92] & (((din_a[91] & din_b[94])))) # (din_a[92] & (!din_b[93] $ (((!din_a[91]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_554  ) + ( Xd_0__inst_mult_7_553  ))
// Xd_0__inst_mult_7_562  = SHARE((din_a[92] & (din_b[93] & (din_a[91] & din_b[94]))))

	.dataa(!din_a[92]),
	.datab(!din_b[93]),
	.datac(!din_a[91]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_553 ),
	.sharein(Xd_0__inst_mult_7_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_560 ),
	.cout(Xd_0__inst_mult_7_561 ),
	.shareout(Xd_0__inst_mult_7_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_167 (
// Equation(s):
// Xd_0__inst_mult_4_568  = SUM(( GND ) + ( Xd_0__inst_mult_4_566  ) + ( Xd_0__inst_mult_4_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_565 ),
	.sharein(Xd_0__inst_mult_4_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_161 (
// Equation(s):
// Xd_0__inst_mult_5_556  = SUM(( GND ) + ( Xd_0__inst_mult_5_550  ) + ( Xd_0__inst_mult_5_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_549 ),
	.sharein(Xd_0__inst_mult_5_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_162 (
// Equation(s):
// Xd_0__inst_mult_5_560  = SUM(( (!din_a[68] & (((din_a[67] & din_b[70])))) # (din_a[68] & (!din_b[69] $ (((!din_a[67]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_554  ) + ( Xd_0__inst_mult_5_553  ))
// Xd_0__inst_mult_5_561  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[70])))) # (din_a[68] & (!din_b[69] $ (((!din_a[67]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_554  ) + ( Xd_0__inst_mult_5_553  ))
// Xd_0__inst_mult_5_562  = SHARE((din_a[68] & (din_b[69] & (din_a[67] & din_b[70]))))

	.dataa(!din_a[68]),
	.datab(!din_b[69]),
	.datac(!din_a[67]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_553 ),
	.sharein(Xd_0__inst_mult_5_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_560 ),
	.cout(Xd_0__inst_mult_5_561 ),
	.shareout(Xd_0__inst_mult_5_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_165 (
// Equation(s):
// Xd_0__inst_mult_2_560  = SUM(( GND ) + ( Xd_0__inst_mult_2_554  ) + ( Xd_0__inst_mult_2_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_553 ),
	.sharein(Xd_0__inst_mult_2_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_166 (
// Equation(s):
// Xd_0__inst_mult_2_564  = SUM(( (!din_a[32] & (((din_a[31] & din_b[34])))) # (din_a[32] & (!din_b[33] $ (((!din_a[31]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_558  ) + ( Xd_0__inst_mult_2_557  ))
// Xd_0__inst_mult_2_565  = CARRY(( (!din_a[32] & (((din_a[31] & din_b[34])))) # (din_a[32] & (!din_b[33] $ (((!din_a[31]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_558  ) + ( Xd_0__inst_mult_2_557  ))
// Xd_0__inst_mult_2_566  = SHARE((din_a[32] & (din_b[33] & (din_a[31] & din_b[34]))))

	.dataa(!din_a[32]),
	.datab(!din_b[33]),
	.datac(!din_a[31]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_557 ),
	.sharein(Xd_0__inst_mult_2_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_564 ),
	.cout(Xd_0__inst_mult_2_565 ),
	.shareout(Xd_0__inst_mult_2_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_161 (
// Equation(s):
// Xd_0__inst_mult_3_556  = SUM(( GND ) + ( Xd_0__inst_mult_3_550  ) + ( Xd_0__inst_mult_3_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_549 ),
	.sharein(Xd_0__inst_mult_3_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_162 (
// Equation(s):
// Xd_0__inst_mult_3_560  = SUM(( (!din_a[44] & (((din_a[43] & din_b[46])))) # (din_a[44] & (!din_b[45] $ (((!din_a[43]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_554  ) + ( Xd_0__inst_mult_3_553  ))
// Xd_0__inst_mult_3_561  = CARRY(( (!din_a[44] & (((din_a[43] & din_b[46])))) # (din_a[44] & (!din_b[45] $ (((!din_a[43]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_554  ) + ( Xd_0__inst_mult_3_553  ))
// Xd_0__inst_mult_3_562  = SHARE((din_a[44] & (din_b[45] & (din_a[43] & din_b[46]))))

	.dataa(!din_a[44]),
	.datab(!din_b[45]),
	.datac(!din_a[43]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_553 ),
	.sharein(Xd_0__inst_mult_3_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_560 ),
	.cout(Xd_0__inst_mult_3_561 ),
	.shareout(Xd_0__inst_mult_3_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_165 (
// Equation(s):
// Xd_0__inst_mult_0_560  = SUM(( GND ) + ( Xd_0__inst_mult_0_554  ) + ( Xd_0__inst_mult_0_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_553 ),
	.sharein(Xd_0__inst_mult_0_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_166 (
// Equation(s):
// Xd_0__inst_mult_0_564  = SUM(( (!din_a[8] & (((din_a[7] & din_b[10])))) # (din_a[8] & (!din_b[9] $ (((!din_a[7]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_558  ) + ( Xd_0__inst_mult_0_557  ))
// Xd_0__inst_mult_0_565  = CARRY(( (!din_a[8] & (((din_a[7] & din_b[10])))) # (din_a[8] & (!din_b[9] $ (((!din_a[7]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_558  ) + ( Xd_0__inst_mult_0_557  ))
// Xd_0__inst_mult_0_566  = SHARE((din_a[8] & (din_b[9] & (din_a[7] & din_b[10]))))

	.dataa(!din_a[8]),
	.datab(!din_b[9]),
	.datac(!din_a[7]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_557 ),
	.sharein(Xd_0__inst_mult_0_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_564 ),
	.cout(Xd_0__inst_mult_0_565 ),
	.shareout(Xd_0__inst_mult_0_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_166 (
// Equation(s):
// Xd_0__inst_mult_1_564  = SUM(( GND ) + ( Xd_0__inst_mult_1_558  ) + ( Xd_0__inst_mult_1_557  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_557 ),
	.sharein(Xd_0__inst_mult_1_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_564 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_167 (
// Equation(s):
// Xd_0__inst_mult_1_568  = SUM(( (!din_a[20] & (((din_a[19] & din_b[22])))) # (din_a[20] & (!din_b[21] $ (((!din_a[19]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_562  ) + ( Xd_0__inst_mult_1_561  ))
// Xd_0__inst_mult_1_569  = CARRY(( (!din_a[20] & (((din_a[19] & din_b[22])))) # (din_a[20] & (!din_b[21] $ (((!din_a[19]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_562  ) + ( Xd_0__inst_mult_1_561  ))
// Xd_0__inst_mult_1_570  = SHARE((din_a[20] & (din_b[21] & (din_a[19] & din_b[22]))))

	.dataa(!din_a[20]),
	.datab(!din_b[21]),
	.datac(!din_a[19]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_561 ),
	.sharein(Xd_0__inst_mult_1_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_568 ),
	.cout(Xd_0__inst_mult_1_569 ),
	.shareout(Xd_0__inst_mult_1_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_167 (
// Equation(s):
// Xd_0__inst_mult_13_568  = SUM(( (din_a[164] & din_b[166]) ) + ( Xd_0__inst_mult_13_566  ) + ( Xd_0__inst_mult_13_565  ))
// Xd_0__inst_mult_13_569  = CARRY(( (din_a[164] & din_b[166]) ) + ( Xd_0__inst_mult_13_566  ) + ( Xd_0__inst_mult_13_565  ))
// Xd_0__inst_mult_13_570  = SHARE(GND)

	.dataa(!din_a[164]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_565 ),
	.sharein(Xd_0__inst_mult_13_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_568 ),
	.cout(Xd_0__inst_mult_13_569 ),
	.shareout(Xd_0__inst_mult_13_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_168 (
// Equation(s):
// Xd_0__inst_mult_14_572  = SUM(( (din_a[176] & din_b[178]) ) + ( Xd_0__inst_mult_14_570  ) + ( Xd_0__inst_mult_14_569  ))
// Xd_0__inst_mult_14_573  = CARRY(( (din_a[176] & din_b[178]) ) + ( Xd_0__inst_mult_14_570  ) + ( Xd_0__inst_mult_14_569  ))
// Xd_0__inst_mult_14_574  = SHARE(GND)

	.dataa(!din_a[176]),
	.datab(!din_b[178]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_569 ),
	.sharein(Xd_0__inst_mult_14_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_572 ),
	.cout(Xd_0__inst_mult_14_573 ),
	.shareout(Xd_0__inst_mult_14_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_163 (
// Equation(s):
// Xd_0__inst_mult_10_564  = SUM(( (din_a[128] & din_b[130]) ) + ( Xd_0__inst_mult_10_562  ) + ( Xd_0__inst_mult_10_561  ))
// Xd_0__inst_mult_10_565  = CARRY(( (din_a[128] & din_b[130]) ) + ( Xd_0__inst_mult_10_562  ) + ( Xd_0__inst_mult_10_561  ))
// Xd_0__inst_mult_10_566  = SHARE(GND)

	.dataa(!din_a[128]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_561 ),
	.sharein(Xd_0__inst_mult_10_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_564 ),
	.cout(Xd_0__inst_mult_10_565 ),
	.shareout(Xd_0__inst_mult_10_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_167 (
// Equation(s):
// Xd_0__inst_mult_11_568  = SUM(( (din_a[140] & din_b[142]) ) + ( Xd_0__inst_mult_11_566  ) + ( Xd_0__inst_mult_11_565  ))
// Xd_0__inst_mult_11_569  = CARRY(( (din_a[140] & din_b[142]) ) + ( Xd_0__inst_mult_11_566  ) + ( Xd_0__inst_mult_11_565  ))
// Xd_0__inst_mult_11_570  = SHARE(GND)

	.dataa(!din_a[140]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_565 ),
	.sharein(Xd_0__inst_mult_11_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_568 ),
	.cout(Xd_0__inst_mult_11_569 ),
	.shareout(Xd_0__inst_mult_11_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_167 (
// Equation(s):
// Xd_0__inst_mult_8_568  = SUM(( (din_a[104] & din_b[106]) ) + ( Xd_0__inst_mult_8_566  ) + ( Xd_0__inst_mult_8_565  ))
// Xd_0__inst_mult_8_569  = CARRY(( (din_a[104] & din_b[106]) ) + ( Xd_0__inst_mult_8_566  ) + ( Xd_0__inst_mult_8_565  ))
// Xd_0__inst_mult_8_570  = SHARE(GND)

	.dataa(!din_a[104]),
	.datab(!din_b[106]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_565 ),
	.sharein(Xd_0__inst_mult_8_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_568 ),
	.cout(Xd_0__inst_mult_8_569 ),
	.shareout(Xd_0__inst_mult_8_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_163 (
// Equation(s):
// Xd_0__inst_mult_9_564  = SUM(( (din_a[116] & din_b[118]) ) + ( Xd_0__inst_mult_9_562  ) + ( Xd_0__inst_mult_9_561  ))
// Xd_0__inst_mult_9_565  = CARRY(( (din_a[116] & din_b[118]) ) + ( Xd_0__inst_mult_9_562  ) + ( Xd_0__inst_mult_9_561  ))
// Xd_0__inst_mult_9_566  = SHARE(GND)

	.dataa(!din_a[116]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_561 ),
	.sharein(Xd_0__inst_mult_9_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_564 ),
	.cout(Xd_0__inst_mult_9_565 ),
	.shareout(Xd_0__inst_mult_9_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_163 (
// Equation(s):
// Xd_0__inst_mult_6_564  = SUM(( (din_a[80] & din_b[82]) ) + ( Xd_0__inst_mult_6_562  ) + ( Xd_0__inst_mult_6_561  ))
// Xd_0__inst_mult_6_565  = CARRY(( (din_a[80] & din_b[82]) ) + ( Xd_0__inst_mult_6_562  ) + ( Xd_0__inst_mult_6_561  ))
// Xd_0__inst_mult_6_566  = SHARE(GND)

	.dataa(!din_a[80]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_561 ),
	.sharein(Xd_0__inst_mult_6_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_564 ),
	.cout(Xd_0__inst_mult_6_565 ),
	.shareout(Xd_0__inst_mult_6_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_163 (
// Equation(s):
// Xd_0__inst_mult_7_564  = SUM(( (din_a[92] & din_b[94]) ) + ( Xd_0__inst_mult_7_562  ) + ( Xd_0__inst_mult_7_561  ))
// Xd_0__inst_mult_7_565  = CARRY(( (din_a[92] & din_b[94]) ) + ( Xd_0__inst_mult_7_562  ) + ( Xd_0__inst_mult_7_561  ))
// Xd_0__inst_mult_7_566  = SHARE(GND)

	.dataa(!din_a[92]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_561 ),
	.sharein(Xd_0__inst_mult_7_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_564 ),
	.cout(Xd_0__inst_mult_7_565 ),
	.shareout(Xd_0__inst_mult_7_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_163 (
// Equation(s):
// Xd_0__inst_mult_5_564  = SUM(( (din_a[68] & din_b[70]) ) + ( Xd_0__inst_mult_5_562  ) + ( Xd_0__inst_mult_5_561  ))
// Xd_0__inst_mult_5_565  = CARRY(( (din_a[68] & din_b[70]) ) + ( Xd_0__inst_mult_5_562  ) + ( Xd_0__inst_mult_5_561  ))
// Xd_0__inst_mult_5_566  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_561 ),
	.sharein(Xd_0__inst_mult_5_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_564 ),
	.cout(Xd_0__inst_mult_5_565 ),
	.shareout(Xd_0__inst_mult_5_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_167 (
// Equation(s):
// Xd_0__inst_mult_2_568  = SUM(( (din_a[32] & din_b[34]) ) + ( Xd_0__inst_mult_2_566  ) + ( Xd_0__inst_mult_2_565  ))
// Xd_0__inst_mult_2_569  = CARRY(( (din_a[32] & din_b[34]) ) + ( Xd_0__inst_mult_2_566  ) + ( Xd_0__inst_mult_2_565  ))
// Xd_0__inst_mult_2_570  = SHARE(GND)

	.dataa(!din_a[32]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_565 ),
	.sharein(Xd_0__inst_mult_2_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_568 ),
	.cout(Xd_0__inst_mult_2_569 ),
	.shareout(Xd_0__inst_mult_2_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_163 (
// Equation(s):
// Xd_0__inst_mult_3_564  = SUM(( (din_a[44] & din_b[46]) ) + ( Xd_0__inst_mult_3_562  ) + ( Xd_0__inst_mult_3_561  ))
// Xd_0__inst_mult_3_565  = CARRY(( (din_a[44] & din_b[46]) ) + ( Xd_0__inst_mult_3_562  ) + ( Xd_0__inst_mult_3_561  ))
// Xd_0__inst_mult_3_566  = SHARE(GND)

	.dataa(!din_a[44]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_561 ),
	.sharein(Xd_0__inst_mult_3_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_564 ),
	.cout(Xd_0__inst_mult_3_565 ),
	.shareout(Xd_0__inst_mult_3_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_167 (
// Equation(s):
// Xd_0__inst_mult_0_568  = SUM(( (din_a[8] & din_b[10]) ) + ( Xd_0__inst_mult_0_566  ) + ( Xd_0__inst_mult_0_565  ))
// Xd_0__inst_mult_0_569  = CARRY(( (din_a[8] & din_b[10]) ) + ( Xd_0__inst_mult_0_566  ) + ( Xd_0__inst_mult_0_565  ))
// Xd_0__inst_mult_0_570  = SHARE(GND)

	.dataa(!din_a[8]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_565 ),
	.sharein(Xd_0__inst_mult_0_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_568 ),
	.cout(Xd_0__inst_mult_0_569 ),
	.shareout(Xd_0__inst_mult_0_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_168 (
// Equation(s):
// Xd_0__inst_mult_1_572  = SUM(( (din_a[20] & din_b[22]) ) + ( Xd_0__inst_mult_1_570  ) + ( Xd_0__inst_mult_1_569  ))
// Xd_0__inst_mult_1_573  = CARRY(( (din_a[20] & din_b[22]) ) + ( Xd_0__inst_mult_1_570  ) + ( Xd_0__inst_mult_1_569  ))
// Xd_0__inst_mult_1_574  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_569 ),
	.sharein(Xd_0__inst_mult_1_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_572 ),
	.cout(Xd_0__inst_mult_1_573 ),
	.shareout(Xd_0__inst_mult_1_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_168 (
// Equation(s):
// Xd_0__inst_mult_13_572  = SUM(( GND ) + ( Xd_0__inst_mult_13_570  ) + ( Xd_0__inst_mult_13_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_569 ),
	.sharein(Xd_0__inst_mult_13_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_169 (
// Equation(s):
// Xd_0__inst_mult_14_576  = SUM(( GND ) + ( Xd_0__inst_mult_14_574  ) + ( Xd_0__inst_mult_14_573  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_573 ),
	.sharein(Xd_0__inst_mult_14_574 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_576 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_164 (
// Equation(s):
// Xd_0__inst_mult_10_568  = SUM(( GND ) + ( Xd_0__inst_mult_10_566  ) + ( Xd_0__inst_mult_10_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_565 ),
	.sharein(Xd_0__inst_mult_10_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_168 (
// Equation(s):
// Xd_0__inst_mult_11_572  = SUM(( GND ) + ( Xd_0__inst_mult_11_570  ) + ( Xd_0__inst_mult_11_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_569 ),
	.sharein(Xd_0__inst_mult_11_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_168 (
// Equation(s):
// Xd_0__inst_mult_8_572  = SUM(( GND ) + ( Xd_0__inst_mult_8_570  ) + ( Xd_0__inst_mult_8_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_569 ),
	.sharein(Xd_0__inst_mult_8_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_164 (
// Equation(s):
// Xd_0__inst_mult_9_568  = SUM(( GND ) + ( Xd_0__inst_mult_9_566  ) + ( Xd_0__inst_mult_9_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_565 ),
	.sharein(Xd_0__inst_mult_9_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_164 (
// Equation(s):
// Xd_0__inst_mult_6_568  = SUM(( GND ) + ( Xd_0__inst_mult_6_566  ) + ( Xd_0__inst_mult_6_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_565 ),
	.sharein(Xd_0__inst_mult_6_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_164 (
// Equation(s):
// Xd_0__inst_mult_7_568  = SUM(( GND ) + ( Xd_0__inst_mult_7_566  ) + ( Xd_0__inst_mult_7_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_565 ),
	.sharein(Xd_0__inst_mult_7_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_164 (
// Equation(s):
// Xd_0__inst_mult_5_568  = SUM(( GND ) + ( Xd_0__inst_mult_5_566  ) + ( Xd_0__inst_mult_5_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_565 ),
	.sharein(Xd_0__inst_mult_5_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_168 (
// Equation(s):
// Xd_0__inst_mult_2_572  = SUM(( GND ) + ( Xd_0__inst_mult_2_570  ) + ( Xd_0__inst_mult_2_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_569 ),
	.sharein(Xd_0__inst_mult_2_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_164 (
// Equation(s):
// Xd_0__inst_mult_3_568  = SUM(( GND ) + ( Xd_0__inst_mult_3_566  ) + ( Xd_0__inst_mult_3_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_565 ),
	.sharein(Xd_0__inst_mult_3_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_168 (
// Equation(s):
// Xd_0__inst_mult_0_572  = SUM(( GND ) + ( Xd_0__inst_mult_0_570  ) + ( Xd_0__inst_mult_0_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_569 ),
	.sharein(Xd_0__inst_mult_0_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_169 (
// Equation(s):
// Xd_0__inst_mult_1_576  = SUM(( GND ) + ( Xd_0__inst_mult_1_574  ) + ( Xd_0__inst_mult_1_573  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_573 ),
	.sharein(Xd_0__inst_mult_1_574 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_576 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_164 (
// Equation(s):
// Xd_0__inst_mult_12_569  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_570  = SHARE((din_a[147] & din_b[145]))

	.dataa(!din_a[147]),
	.datab(!din_b[145]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_569 ),
	.shareout(Xd_0__inst_mult_12_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_169 (
// Equation(s):
// Xd_0__inst_mult_13_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_578  = SHARE((din_a[159] & din_b[157]))

	.dataa(!din_a[159]),
	.datab(!din_b[157]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_577 ),
	.shareout(Xd_0__inst_mult_13_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_165 (
// Equation(s):
// Xd_0__inst_mult_10_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_574  = SHARE((din_a[123] & din_b[121]))

	.dataa(!din_a[123]),
	.datab(!din_b[121]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_573 ),
	.shareout(Xd_0__inst_mult_10_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_169 (
// Equation(s):
// Xd_0__inst_mult_11_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_578  = SHARE((din_a[135] & din_b[133]))

	.dataa(!din_a[135]),
	.datab(!din_b[133]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_577 ),
	.shareout(Xd_0__inst_mult_11_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_169 (
// Equation(s):
// Xd_0__inst_mult_8_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_578  = SHARE((din_a[99] & din_b[97]))

	.dataa(!din_a[99]),
	.datab(!din_b[97]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_577 ),
	.shareout(Xd_0__inst_mult_8_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_165 (
// Equation(s):
// Xd_0__inst_mult_9_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_574  = SHARE((din_a[111] & din_b[109]))

	.dataa(!din_a[111]),
	.datab(!din_b[109]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_573 ),
	.shareout(Xd_0__inst_mult_9_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_165 (
// Equation(s):
// Xd_0__inst_mult_6_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_574  = SHARE((din_a[75] & din_b[73]))

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_573 ),
	.shareout(Xd_0__inst_mult_6_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_165 (
// Equation(s):
// Xd_0__inst_mult_7_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_574  = SHARE((din_a[87] & din_b[85]))

	.dataa(!din_a[87]),
	.datab(!din_b[85]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_573 ),
	.shareout(Xd_0__inst_mult_7_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_168 (
// Equation(s):
// Xd_0__inst_mult_4_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_574  = SHARE((din_a[51] & din_b[49]))

	.dataa(!din_a[51]),
	.datab(!din_b[49]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_573 ),
	.shareout(Xd_0__inst_mult_4_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_165 (
// Equation(s):
// Xd_0__inst_mult_5_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_574  = SHARE((din_a[63] & din_b[61]))

	.dataa(!din_a[63]),
	.datab(!din_b[61]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_573 ),
	.shareout(Xd_0__inst_mult_5_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_169 (
// Equation(s):
// Xd_0__inst_mult_2_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_578  = SHARE((din_a[27] & din_b[25]))

	.dataa(!din_a[27]),
	.datab(!din_b[25]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_577 ),
	.shareout(Xd_0__inst_mult_2_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_165 (
// Equation(s):
// Xd_0__inst_mult_3_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_574  = SHARE((din_a[39] & din_b[37]))

	.dataa(!din_a[39]),
	.datab(!din_b[37]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_573 ),
	.shareout(Xd_0__inst_mult_3_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_169 (
// Equation(s):
// Xd_0__inst_mult_0_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_578  = SHARE((din_a[3] & din_b[1]))

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_577 ),
	.shareout(Xd_0__inst_mult_0_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_165 (
// Equation(s):
// Xd_0__inst_mult_12_573  = CARRY(( (din_a[146] & din_b[151]) ) + ( Xd_0__inst_mult_12_582  ) + ( Xd_0__inst_mult_12_581  ))
// Xd_0__inst_mult_12_574  = SHARE((din_a[145] & din_b[152]))

	.dataa(!din_a[146]),
	.datab(!din_b[151]),
	.datac(!din_a[145]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_581 ),
	.sharein(Xd_0__inst_mult_12_582 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_573 ),
	.shareout(Xd_0__inst_mult_12_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_170 (
// Equation(s):
// Xd_0__inst_mult_13_581  = CARRY(( (din_a[158] & din_b[163]) ) + ( Xd_0__inst_mult_13_550  ) + ( Xd_0__inst_mult_13_549  ))
// Xd_0__inst_mult_13_582  = SHARE((din_a[157] & din_b[164]))

	.dataa(!din_a[158]),
	.datab(!din_b[163]),
	.datac(!din_a[157]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_549 ),
	.sharein(Xd_0__inst_mult_13_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_581 ),
	.shareout(Xd_0__inst_mult_13_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_170 (
// Equation(s):
// Xd_0__inst_mult_14_581  = CARRY(( (din_a[170] & din_b[175]) ) + ( Xd_0__inst_mult_14_542  ) + ( Xd_0__inst_mult_14_541  ))
// Xd_0__inst_mult_14_582  = SHARE((din_a[169] & din_b[176]))

	.dataa(!din_a[170]),
	.datab(!din_b[175]),
	.datac(!din_a[169]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_541 ),
	.sharein(Xd_0__inst_mult_14_542 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_581 ),
	.shareout(Xd_0__inst_mult_14_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_169 (
// Equation(s):
// Xd_0__inst_mult_15_577  = CARRY(( (din_a[182] & din_b[187]) ) + ( Xd_0__inst_mult_15_586  ) + ( Xd_0__inst_mult_15_585  ))
// Xd_0__inst_mult_15_578  = SHARE((din_a[181] & din_b[188]))

	.dataa(!din_a[182]),
	.datab(!din_b[187]),
	.datac(!din_a[181]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_585 ),
	.sharein(Xd_0__inst_mult_15_586 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_577 ),
	.shareout(Xd_0__inst_mult_15_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_166 (
// Equation(s):
// Xd_0__inst_mult_10_577  = CARRY(( (din_a[122] & din_b[127]) ) + ( Xd_0__inst_mult_10_546  ) + ( Xd_0__inst_mult_10_545  ))
// Xd_0__inst_mult_10_578  = SHARE((din_a[121] & din_b[128]))

	.dataa(!din_a[122]),
	.datab(!din_b[127]),
	.datac(!din_a[121]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_545 ),
	.sharein(Xd_0__inst_mult_10_546 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_577 ),
	.shareout(Xd_0__inst_mult_10_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_170 (
// Equation(s):
// Xd_0__inst_mult_11_581  = CARRY(( (din_a[134] & din_b[139]) ) + ( Xd_0__inst_mult_11_550  ) + ( Xd_0__inst_mult_11_549  ))
// Xd_0__inst_mult_11_582  = SHARE((din_a[133] & din_b[140]))

	.dataa(!din_a[134]),
	.datab(!din_b[139]),
	.datac(!din_a[133]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_549 ),
	.sharein(Xd_0__inst_mult_11_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_581 ),
	.shareout(Xd_0__inst_mult_11_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_170 (
// Equation(s):
// Xd_0__inst_mult_8_581  = CARRY(( (din_a[98] & din_b[103]) ) + ( Xd_0__inst_mult_8_550  ) + ( Xd_0__inst_mult_8_549  ))
// Xd_0__inst_mult_8_582  = SHARE((din_a[97] & din_b[104]))

	.dataa(!din_a[98]),
	.datab(!din_b[103]),
	.datac(!din_a[97]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_549 ),
	.sharein(Xd_0__inst_mult_8_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_581 ),
	.shareout(Xd_0__inst_mult_8_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_166 (
// Equation(s):
// Xd_0__inst_mult_9_577  = CARRY(( (din_a[110] & din_b[115]) ) + ( Xd_0__inst_mult_9_546  ) + ( Xd_0__inst_mult_9_545  ))
// Xd_0__inst_mult_9_578  = SHARE((din_a[109] & din_b[116]))

	.dataa(!din_a[110]),
	.datab(!din_b[115]),
	.datac(!din_a[109]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_545 ),
	.sharein(Xd_0__inst_mult_9_546 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_577 ),
	.shareout(Xd_0__inst_mult_9_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_166 (
// Equation(s):
// Xd_0__inst_mult_6_577  = CARRY(( (din_a[74] & din_b[79]) ) + ( Xd_0__inst_mult_6_546  ) + ( Xd_0__inst_mult_6_545  ))
// Xd_0__inst_mult_6_578  = SHARE((din_a[73] & din_b[80]))

	.dataa(!din_a[74]),
	.datab(!din_b[79]),
	.datac(!din_a[73]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_545 ),
	.sharein(Xd_0__inst_mult_6_546 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_577 ),
	.shareout(Xd_0__inst_mult_6_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_166 (
// Equation(s):
// Xd_0__inst_mult_7_577  = CARRY(( (din_a[86] & din_b[91]) ) + ( Xd_0__inst_mult_7_546  ) + ( Xd_0__inst_mult_7_545  ))
// Xd_0__inst_mult_7_578  = SHARE((din_a[85] & din_b[92]))

	.dataa(!din_a[86]),
	.datab(!din_b[91]),
	.datac(!din_a[85]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_545 ),
	.sharein(Xd_0__inst_mult_7_546 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_577 ),
	.shareout(Xd_0__inst_mult_7_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_169 (
// Equation(s):
// Xd_0__inst_mult_4_577  = CARRY(( (din_a[50] & din_b[55]) ) + ( Xd_0__inst_mult_4_586  ) + ( Xd_0__inst_mult_4_585  ))
// Xd_0__inst_mult_4_578  = SHARE((din_a[49] & din_b[56]))

	.dataa(!din_a[50]),
	.datab(!din_b[55]),
	.datac(!din_a[49]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_585 ),
	.sharein(Xd_0__inst_mult_4_586 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_577 ),
	.shareout(Xd_0__inst_mult_4_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_166 (
// Equation(s):
// Xd_0__inst_mult_5_577  = CARRY(( (din_a[62] & din_b[67]) ) + ( Xd_0__inst_mult_5_538  ) + ( Xd_0__inst_mult_5_537  ))
// Xd_0__inst_mult_5_578  = SHARE((din_a[61] & din_b[68]))

	.dataa(!din_a[62]),
	.datab(!din_b[67]),
	.datac(!din_a[61]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_537 ),
	.sharein(Xd_0__inst_mult_5_538 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_577 ),
	.shareout(Xd_0__inst_mult_5_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_170 (
// Equation(s):
// Xd_0__inst_mult_2_581  = CARRY(( (din_a[26] & din_b[31]) ) + ( Xd_0__inst_mult_2_542  ) + ( Xd_0__inst_mult_2_541  ))
// Xd_0__inst_mult_2_582  = SHARE((din_a[25] & din_b[32]))

	.dataa(!din_a[26]),
	.datab(!din_b[31]),
	.datac(!din_a[25]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_541 ),
	.sharein(Xd_0__inst_mult_2_542 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_581 ),
	.shareout(Xd_0__inst_mult_2_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_166 (
// Equation(s):
// Xd_0__inst_mult_3_577  = CARRY(( (din_a[38] & din_b[43]) ) + ( Xd_0__inst_mult_3_538  ) + ( Xd_0__inst_mult_3_537  ))
// Xd_0__inst_mult_3_578  = SHARE((din_a[37] & din_b[44]))

	.dataa(!din_a[38]),
	.datab(!din_b[43]),
	.datac(!din_a[37]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_537 ),
	.sharein(Xd_0__inst_mult_3_538 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_577 ),
	.shareout(Xd_0__inst_mult_3_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_170 (
// Equation(s):
// Xd_0__inst_mult_0_581  = CARRY(( (din_a[2] & din_b[7]) ) + ( Xd_0__inst_mult_0_542  ) + ( Xd_0__inst_mult_0_541  ))
// Xd_0__inst_mult_0_582  = SHARE((din_a[1] & din_b[8]))

	.dataa(!din_a[2]),
	.datab(!din_b[7]),
	.datac(!din_a[1]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_541 ),
	.sharein(Xd_0__inst_mult_0_542 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_581 ),
	.shareout(Xd_0__inst_mult_0_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_170 (
// Equation(s):
// Xd_0__inst_mult_1_581  = CARRY(( (din_a[14] & din_b[19]) ) + ( Xd_0__inst_mult_1_546  ) + ( Xd_0__inst_mult_1_545  ))
// Xd_0__inst_mult_1_582  = SHARE((din_a[13] & din_b[20]))

	.dataa(!din_a[14]),
	.datab(!din_b[19]),
	.datac(!din_a[13]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_545 ),
	.sharein(Xd_0__inst_mult_1_546 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_581 ),
	.shareout(Xd_0__inst_mult_1_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_166 (
// Equation(s):
// Xd_0__inst_mult_12_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_578  = SHARE((din_a[148] & din_b[150]))

	.dataa(!din_a[148]),
	.datab(!din_b[150]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_577 ),
	.shareout(Xd_0__inst_mult_12_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_171 (
// Equation(s):
// Xd_0__inst_mult_13_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_586  = SHARE((din_a[160] & din_b[162]))

	.dataa(!din_a[160]),
	.datab(!din_b[162]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_585 ),
	.shareout(Xd_0__inst_mult_13_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_171 (
// Equation(s):
// Xd_0__inst_mult_14_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_586  = SHARE((din_a[172] & din_b[174]))

	.dataa(!din_a[172]),
	.datab(!din_b[174]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_585 ),
	.shareout(Xd_0__inst_mult_14_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_170 (
// Equation(s):
// Xd_0__inst_mult_15_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_582  = SHARE((din_a[184] & din_b[186]))

	.dataa(!din_a[184]),
	.datab(!din_b[186]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_581 ),
	.shareout(Xd_0__inst_mult_15_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_167 (
// Equation(s):
// Xd_0__inst_mult_10_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_582  = SHARE((din_a[124] & din_b[126]))

	.dataa(!din_a[124]),
	.datab(!din_b[126]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_581 ),
	.shareout(Xd_0__inst_mult_10_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_171 (
// Equation(s):
// Xd_0__inst_mult_11_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_586  = SHARE((din_a[136] & din_b[138]))

	.dataa(!din_a[136]),
	.datab(!din_b[138]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_585 ),
	.shareout(Xd_0__inst_mult_11_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_171 (
// Equation(s):
// Xd_0__inst_mult_8_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_586  = SHARE((din_a[100] & din_b[102]))

	.dataa(!din_a[100]),
	.datab(!din_b[102]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_585 ),
	.shareout(Xd_0__inst_mult_8_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_167 (
// Equation(s):
// Xd_0__inst_mult_9_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_582  = SHARE((din_a[112] & din_b[114]))

	.dataa(!din_a[112]),
	.datab(!din_b[114]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_581 ),
	.shareout(Xd_0__inst_mult_9_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_167 (
// Equation(s):
// Xd_0__inst_mult_6_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_582  = SHARE((din_a[76] & din_b[78]))

	.dataa(!din_a[76]),
	.datab(!din_b[78]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_581 ),
	.shareout(Xd_0__inst_mult_6_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_167 (
// Equation(s):
// Xd_0__inst_mult_7_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_582  = SHARE((din_a[88] & din_b[90]))

	.dataa(!din_a[88]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_581 ),
	.shareout(Xd_0__inst_mult_7_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_170 (
// Equation(s):
// Xd_0__inst_mult_4_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_582  = SHARE((din_a[52] & din_b[54]))

	.dataa(!din_a[52]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_581 ),
	.shareout(Xd_0__inst_mult_4_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_167 (
// Equation(s):
// Xd_0__inst_mult_5_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_582  = SHARE((din_a[64] & din_b[66]))

	.dataa(!din_a[64]),
	.datab(!din_b[66]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_581 ),
	.shareout(Xd_0__inst_mult_5_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_171 (
// Equation(s):
// Xd_0__inst_mult_2_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_586  = SHARE((din_a[28] & din_b[30]))

	.dataa(!din_a[28]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_585 ),
	.shareout(Xd_0__inst_mult_2_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_167 (
// Equation(s):
// Xd_0__inst_mult_3_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_582  = SHARE((din_a[40] & din_b[42]))

	.dataa(!din_a[40]),
	.datab(!din_b[42]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_581 ),
	.shareout(Xd_0__inst_mult_3_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_171 (
// Equation(s):
// Xd_0__inst_mult_0_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_586  = SHARE((din_a[4] & din_b[6]))

	.dataa(!din_a[4]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_585 ),
	.shareout(Xd_0__inst_mult_0_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_171 (
// Equation(s):
// Xd_0__inst_mult_1_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_586  = SHARE((din_a[16] & din_b[18]))

	.dataa(!din_a[16]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_585 ),
	.shareout(Xd_0__inst_mult_1_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_167 (
// Equation(s):
// Xd_0__inst_mult_12_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_582  = SHARE((din_a[146] & din_b[151]))

	.dataa(!din_a[146]),
	.datab(!din_b[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_581 ),
	.shareout(Xd_0__inst_mult_12_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_171 (
// Equation(s):
// Xd_0__inst_mult_15_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_586  = SHARE((din_a[182] & din_b[187]))

	.dataa(!din_a[182]),
	.datab(!din_b[187]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_585 ),
	.shareout(Xd_0__inst_mult_15_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_171 (
// Equation(s):
// Xd_0__inst_mult_4_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_586  = SHARE((din_a[50] & din_b[55]))

	.dataa(!din_a[50]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_585 ),
	.shareout(Xd_0__inst_mult_4_586 ));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [18]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [19]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [20]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [21]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [22]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [23]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [24]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [25]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_26_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_rtl_105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [26]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__25__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__24__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__24__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__25__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__25__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_12_ (
	.clk(clk),
	.d(Xd_0__inst_i29_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_13_ (
	.clk(clk),
	.d(Xd_0__inst_i29_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_14_ (
	.clk(clk),
	.d(Xd_0__inst_i29_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_15_ (
	.clk(clk),
	.d(Xd_0__inst_i29_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_10_ (
	.clk(clk),
	.d(Xd_0__inst_i29_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_11_ (
	.clk(clk),
	.d(Xd_0__inst_i29_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_8_ (
	.clk(clk),
	.d(Xd_0__inst_i29_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_9_ (
	.clk(clk),
	.d(Xd_0__inst_i29_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_6_ (
	.clk(clk),
	.d(Xd_0__inst_i29_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_7_ (
	.clk(clk),
	.d(Xd_0__inst_i29_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_4_ (
	.clk(clk),
	.d(Xd_0__inst_i29_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_5_ (
	.clk(clk),
	.d(Xd_0__inst_i29_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_2_ (
	.clk(clk),
	.d(Xd_0__inst_i29_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_3_ (
	.clk(clk),
	.d(Xd_0__inst_i29_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_0_ (
	.clk(clk),
	.d(Xd_0__inst_i29_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_1_ (
	.clk(clk),
	.d(Xd_0__inst_i29_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_22 (
	.clk(clk),
	.d(din_a[154]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_23 (
	.clk(clk),
	.d(din_b[149]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_22 (
	.clk(clk),
	.d(din_a[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_23 (
	.clk(clk),
	.d(din_b[161]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_22 (
	.clk(clk),
	.d(din_a[178]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_23 (
	.clk(clk),
	.d(din_b[173]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_388 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_22 (
	.clk(clk),
	.d(din_a[190]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_23 (
	.clk(clk),
	.d(din_b[185]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_22 (
	.clk(clk),
	.d(din_a[130]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_23 (
	.clk(clk),
	.d(din_b[125]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_22 (
	.clk(clk),
	.d(din_a[142]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_23 (
	.clk(clk),
	.d(din_b[137]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_22 (
	.clk(clk),
	.d(din_a[106]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_23 (
	.clk(clk),
	.d(din_b[101]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_22 (
	.clk(clk),
	.d(din_a[118]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_23 (
	.clk(clk),
	.d(din_b[113]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_22 (
	.clk(clk),
	.d(din_a[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_23 (
	.clk(clk),
	.d(din_b[77]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_22 (
	.clk(clk),
	.d(din_a[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_23 (
	.clk(clk),
	.d(din_b[89]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_388 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_22 (
	.clk(clk),
	.d(din_a[58]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_23 (
	.clk(clk),
	.d(din_b[53]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_22 (
	.clk(clk),
	.d(din_a[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_23 (
	.clk(clk),
	.d(din_b[65]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_22 (
	.clk(clk),
	.d(din_a[34]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_23 (
	.clk(clk),
	.d(din_b[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_22 (
	.clk(clk),
	.d(din_a[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_23 (
	.clk(clk),
	.d(din_b[41]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_22 (
	.clk(clk),
	.d(din_a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_23 (
	.clk(clk),
	.d(din_b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_22 (
	.clk(clk),
	.d(din_a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_23 (
	.clk(clk),
	.d(din_b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_388 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_392 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_392 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_392 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_388 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_396 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_396 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_396 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_392 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_400 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_400 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_400 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_396 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_63_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_400 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_408 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_408 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_33_q ),
	.prn(vcc));

assign dout[0] = Xd_0__inst_inst_inst_dout [0];

assign dout[1] = Xd_0__inst_inst_inst_dout [1];

assign dout[2] = Xd_0__inst_inst_inst_dout [2];

assign dout[3] = Xd_0__inst_inst_inst_dout [3];

assign dout[4] = Xd_0__inst_inst_inst_dout [4];

assign dout[5] = Xd_0__inst_inst_inst_dout [5];

assign dout[6] = Xd_0__inst_inst_inst_dout [6];

assign dout[7] = Xd_0__inst_inst_inst_dout [7];

assign dout[8] = Xd_0__inst_inst_inst_dout [8];

assign dout[9] = Xd_0__inst_inst_inst_dout [9];

assign dout[10] = Xd_0__inst_inst_inst_dout [10];

assign dout[11] = Xd_0__inst_inst_inst_dout [11];

assign dout[12] = Xd_0__inst_inst_inst_dout [12];

assign dout[13] = Xd_0__inst_inst_inst_dout [13];

assign dout[14] = Xd_0__inst_inst_inst_dout [14];

assign dout[15] = Xd_0__inst_inst_inst_dout [15];

assign dout[16] = Xd_0__inst_inst_inst_dout [16];

assign dout[17] = Xd_0__inst_inst_inst_dout [17];

assign dout[18] = Xd_0__inst_inst_inst_dout [18];

assign dout[19] = Xd_0__inst_inst_inst_dout [19];

assign dout[20] = Xd_0__inst_inst_inst_dout [20];

assign dout[21] = Xd_0__inst_inst_inst_dout [21];

assign dout[22] = Xd_0__inst_inst_inst_dout [22];

assign dout[23] = Xd_0__inst_inst_inst_dout [23];

assign dout[24] = Xd_0__inst_inst_inst_dout [24];

assign dout[25] = Xd_0__inst_inst_inst_dout [25];

assign dout[26] = Xd_0__inst_inst_inst_dout [26];

endmodule
