// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Internal Build 259 12/02/2018 SJ Pro Edition"

// DATE "12/08/2018 22:50:54"

// 
// Device: Altera 1SG280LU2F50E2VG Package FBGA2397
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module pe_dot_alm_s10_8x8x32 (
	dout,
	clk,
	din_a,
	din_b);
output 	[19:0] dout;
input 	clk;
input 	[255:0] din_a;
input 	[255:0] din_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire Xd_0__inst_inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_inst_add_0_6_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_inst_add_0_11_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_12 ;
wire Xd_0__inst_inst_inst_inst_add_0_16_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_17 ;
wire Xd_0__inst_inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_inst_add_0_26_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_inst_add_0_31_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_32 ;
wire Xd_0__inst_inst_inst_inst_add_0_36_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_37 ;
wire Xd_0__inst_inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_inst_add_0_46_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_inst_add_0_51_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_52 ;
wire Xd_0__inst_inst_inst_inst_add_0_56_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_57 ;
wire Xd_0__inst_inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_inst_add_0_66_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_67 ;
wire Xd_0__inst_inst_inst_inst_add_0_71_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_72 ;
wire Xd_0__inst_inst_inst_inst_add_0_76_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_77 ;
wire Xd_0__inst_inst_inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_82 ;
wire Xd_0__inst_inst_inst_inst_add_0_86_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_87 ;
wire Xd_0__inst_inst_inst_inst_add_0_91_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_92 ;
wire Xd_0__inst_inst_inst_inst_add_0_96_sumout ;
wire Xd_0__inst_inst_inst_add_1_1_sumout ;
wire Xd_0__inst_inst_inst_add_1_2 ;
wire Xd_0__inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_add_1_6_sumout ;
wire Xd_0__inst_inst_inst_add_1_7 ;
wire Xd_0__inst_inst_inst_add_0_6_sumout ;
wire Xd_0__inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_add_1_11_sumout ;
wire Xd_0__inst_inst_inst_add_1_12 ;
wire Xd_0__inst_inst_inst_add_0_11_sumout ;
wire Xd_0__inst_inst_inst_add_0_12 ;
wire Xd_0__inst_inst_inst_add_1_16_sumout ;
wire Xd_0__inst_inst_inst_add_1_17 ;
wire Xd_0__inst_inst_inst_add_0_16_sumout ;
wire Xd_0__inst_inst_inst_add_0_17 ;
wire Xd_0__inst_inst_inst_add_1_21_sumout ;
wire Xd_0__inst_inst_inst_add_1_22 ;
wire Xd_0__inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_add_1_26_sumout ;
wire Xd_0__inst_inst_inst_add_1_27 ;
wire Xd_0__inst_inst_inst_add_0_26_sumout ;
wire Xd_0__inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_add_1_31_sumout ;
wire Xd_0__inst_inst_inst_add_1_32 ;
wire Xd_0__inst_inst_inst_add_0_31_sumout ;
wire Xd_0__inst_inst_inst_add_0_32 ;
wire Xd_0__inst_inst_inst_add_1_36_sumout ;
wire Xd_0__inst_inst_inst_add_1_37 ;
wire Xd_0__inst_inst_inst_add_0_36_sumout ;
wire Xd_0__inst_inst_inst_add_0_37 ;
wire Xd_0__inst_inst_inst_add_1_41_sumout ;
wire Xd_0__inst_inst_inst_add_1_42 ;
wire Xd_0__inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_add_1_46_sumout ;
wire Xd_0__inst_inst_inst_add_1_47 ;
wire Xd_0__inst_inst_inst_add_0_46_sumout ;
wire Xd_0__inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_add_1_51_sumout ;
wire Xd_0__inst_inst_inst_add_1_52 ;
wire Xd_0__inst_inst_inst_add_0_51_sumout ;
wire Xd_0__inst_inst_inst_add_0_52 ;
wire Xd_0__inst_inst_inst_add_1_56_sumout ;
wire Xd_0__inst_inst_inst_add_1_57 ;
wire Xd_0__inst_inst_inst_add_0_56_sumout ;
wire Xd_0__inst_inst_inst_add_0_57 ;
wire Xd_0__inst_inst_inst_add_1_61_sumout ;
wire Xd_0__inst_inst_inst_add_1_62 ;
wire Xd_0__inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_add_1_66_sumout ;
wire Xd_0__inst_inst_inst_add_1_67 ;
wire Xd_0__inst_inst_inst_add_0_66_sumout ;
wire Xd_0__inst_inst_inst_add_0_67 ;
wire Xd_0__inst_inst_inst_add_1_71_sumout ;
wire Xd_0__inst_inst_inst_add_1_72 ;
wire Xd_0__inst_inst_inst_add_0_71_sumout ;
wire Xd_0__inst_inst_inst_add_0_72 ;
wire Xd_0__inst_inst_inst_add_1_76_sumout ;
wire Xd_0__inst_inst_inst_add_1_77 ;
wire Xd_0__inst_inst_inst_add_0_76_sumout ;
wire Xd_0__inst_inst_inst_add_0_77 ;
wire Xd_0__inst_inst_inst_add_1_81_sumout ;
wire Xd_0__inst_inst_inst_add_1_82 ;
wire Xd_0__inst_inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_inst_add_0_82 ;
wire Xd_0__inst_inst_inst_add_1_86_sumout ;
wire Xd_0__inst_inst_inst_add_1_87 ;
wire Xd_0__inst_inst_inst_add_0_86_sumout ;
wire Xd_0__inst_inst_inst_add_0_87 ;
wire Xd_0__inst_inst_inst_add_1_91_sumout ;
wire Xd_0__inst_inst_inst_add_0_91_sumout ;
wire Xd_0__inst_mult_12_23_sumout ;
wire Xd_0__inst_mult_12_24 ;
wire Xd_0__inst_mult_13_23_sumout ;
wire Xd_0__inst_mult_13_24 ;
wire Xd_0__inst_inst_add_3_1_sumout ;
wire Xd_0__inst_inst_add_3_2 ;
wire Xd_0__inst_inst_add_2_1_sumout ;
wire Xd_0__inst_inst_add_2_2 ;
wire Xd_0__inst_inst_add_1_1_sumout ;
wire Xd_0__inst_inst_add_1_2 ;
wire Xd_0__inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_add_0_2 ;
wire Xd_0__inst_inst_add_3_6_sumout ;
wire Xd_0__inst_inst_add_3_7 ;
wire Xd_0__inst_inst_add_2_6_sumout ;
wire Xd_0__inst_inst_add_2_7 ;
wire Xd_0__inst_inst_add_1_6_sumout ;
wire Xd_0__inst_inst_add_1_7 ;
wire Xd_0__inst_inst_add_0_6_sumout ;
wire Xd_0__inst_inst_add_0_7 ;
wire Xd_0__inst_inst_add_3_11_sumout ;
wire Xd_0__inst_inst_add_3_12 ;
wire Xd_0__inst_inst_add_2_11_sumout ;
wire Xd_0__inst_inst_add_2_12 ;
wire Xd_0__inst_inst_add_1_11_sumout ;
wire Xd_0__inst_inst_add_1_12 ;
wire Xd_0__inst_inst_add_0_11_sumout ;
wire Xd_0__inst_inst_add_0_12 ;
wire Xd_0__inst_inst_add_3_16_sumout ;
wire Xd_0__inst_inst_add_3_17 ;
wire Xd_0__inst_inst_add_2_16_sumout ;
wire Xd_0__inst_inst_add_2_17 ;
wire Xd_0__inst_inst_add_1_16_sumout ;
wire Xd_0__inst_inst_add_1_17 ;
wire Xd_0__inst_inst_add_0_16_sumout ;
wire Xd_0__inst_inst_add_0_17 ;
wire Xd_0__inst_inst_add_3_21_sumout ;
wire Xd_0__inst_inst_add_3_22 ;
wire Xd_0__inst_inst_add_2_21_sumout ;
wire Xd_0__inst_inst_add_2_22 ;
wire Xd_0__inst_inst_add_1_21_sumout ;
wire Xd_0__inst_inst_add_1_22 ;
wire Xd_0__inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_add_0_22 ;
wire Xd_0__inst_inst_add_3_26_sumout ;
wire Xd_0__inst_inst_add_3_27 ;
wire Xd_0__inst_inst_add_2_26_sumout ;
wire Xd_0__inst_inst_add_2_27 ;
wire Xd_0__inst_inst_add_1_26_sumout ;
wire Xd_0__inst_inst_add_1_27 ;
wire Xd_0__inst_inst_add_0_26_sumout ;
wire Xd_0__inst_inst_add_0_27 ;
wire Xd_0__inst_inst_add_3_31_sumout ;
wire Xd_0__inst_inst_add_3_32 ;
wire Xd_0__inst_inst_add_2_31_sumout ;
wire Xd_0__inst_inst_add_2_32 ;
wire Xd_0__inst_inst_add_1_31_sumout ;
wire Xd_0__inst_inst_add_1_32 ;
wire Xd_0__inst_inst_add_0_31_sumout ;
wire Xd_0__inst_inst_add_0_32 ;
wire Xd_0__inst_inst_add_3_36_sumout ;
wire Xd_0__inst_inst_add_3_37 ;
wire Xd_0__inst_inst_add_2_36_sumout ;
wire Xd_0__inst_inst_add_2_37 ;
wire Xd_0__inst_inst_add_1_36_sumout ;
wire Xd_0__inst_inst_add_1_37 ;
wire Xd_0__inst_inst_add_0_36_sumout ;
wire Xd_0__inst_inst_add_0_37 ;
wire Xd_0__inst_inst_add_3_41_sumout ;
wire Xd_0__inst_inst_add_3_42 ;
wire Xd_0__inst_inst_add_2_41_sumout ;
wire Xd_0__inst_inst_add_2_42 ;
wire Xd_0__inst_inst_add_1_41_sumout ;
wire Xd_0__inst_inst_add_1_42 ;
wire Xd_0__inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_add_0_42 ;
wire Xd_0__inst_inst_add_3_46_sumout ;
wire Xd_0__inst_inst_add_3_47 ;
wire Xd_0__inst_inst_add_2_46_sumout ;
wire Xd_0__inst_inst_add_2_47 ;
wire Xd_0__inst_inst_add_1_46_sumout ;
wire Xd_0__inst_inst_add_1_47 ;
wire Xd_0__inst_inst_add_0_46_sumout ;
wire Xd_0__inst_inst_add_0_47 ;
wire Xd_0__inst_inst_add_3_51_sumout ;
wire Xd_0__inst_inst_add_3_52 ;
wire Xd_0__inst_inst_add_2_51_sumout ;
wire Xd_0__inst_inst_add_2_52 ;
wire Xd_0__inst_inst_add_1_51_sumout ;
wire Xd_0__inst_inst_add_1_52 ;
wire Xd_0__inst_inst_add_0_51_sumout ;
wire Xd_0__inst_inst_add_0_52 ;
wire Xd_0__inst_inst_add_3_56_sumout ;
wire Xd_0__inst_inst_add_3_57 ;
wire Xd_0__inst_inst_add_2_56_sumout ;
wire Xd_0__inst_inst_add_2_57 ;
wire Xd_0__inst_inst_add_1_56_sumout ;
wire Xd_0__inst_inst_add_1_57 ;
wire Xd_0__inst_inst_add_0_56_sumout ;
wire Xd_0__inst_inst_add_0_57 ;
wire Xd_0__inst_inst_add_3_61_sumout ;
wire Xd_0__inst_inst_add_3_62 ;
wire Xd_0__inst_inst_add_2_61_sumout ;
wire Xd_0__inst_inst_add_2_62 ;
wire Xd_0__inst_inst_add_1_61_sumout ;
wire Xd_0__inst_inst_add_1_62 ;
wire Xd_0__inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_add_0_62 ;
wire Xd_0__inst_inst_add_3_66_sumout ;
wire Xd_0__inst_inst_add_3_67 ;
wire Xd_0__inst_inst_add_2_66_sumout ;
wire Xd_0__inst_inst_add_2_67 ;
wire Xd_0__inst_inst_add_1_66_sumout ;
wire Xd_0__inst_inst_add_1_67 ;
wire Xd_0__inst_inst_add_0_66_sumout ;
wire Xd_0__inst_inst_add_0_67 ;
wire Xd_0__inst_inst_add_3_71_sumout ;
wire Xd_0__inst_inst_add_3_72 ;
wire Xd_0__inst_inst_add_2_71_sumout ;
wire Xd_0__inst_inst_add_2_72 ;
wire Xd_0__inst_inst_add_1_71_sumout ;
wire Xd_0__inst_inst_add_1_72 ;
wire Xd_0__inst_inst_add_0_71_sumout ;
wire Xd_0__inst_inst_add_0_72 ;
wire Xd_0__inst_inst_add_3_76_sumout ;
wire Xd_0__inst_inst_add_3_77 ;
wire Xd_0__inst_inst_add_2_76_sumout ;
wire Xd_0__inst_inst_add_2_77 ;
wire Xd_0__inst_inst_add_1_76_sumout ;
wire Xd_0__inst_inst_add_1_77 ;
wire Xd_0__inst_inst_add_0_76_sumout ;
wire Xd_0__inst_inst_add_0_77 ;
wire Xd_0__inst_inst_add_3_81_sumout ;
wire Xd_0__inst_inst_add_3_82 ;
wire Xd_0__inst_inst_add_2_81_sumout ;
wire Xd_0__inst_inst_add_2_82 ;
wire Xd_0__inst_inst_add_1_81_sumout ;
wire Xd_0__inst_inst_add_1_82 ;
wire Xd_0__inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_add_0_82 ;
wire Xd_0__inst_inst_add_3_86_sumout ;
wire Xd_0__inst_inst_add_2_86_sumout ;
wire Xd_0__inst_inst_add_1_86_sumout ;
wire Xd_0__inst_inst_add_0_86_sumout ;
wire Xd_0__inst_mult_11_23_sumout ;
wire Xd_0__inst_mult_11_24 ;
wire Xd_0__inst_mult_22_23_sumout ;
wire Xd_0__inst_mult_22_24 ;
wire Xd_0__inst_mult_24_23_sumout ;
wire Xd_0__inst_mult_24_24 ;
wire Xd_0__inst_mult_26_23_sumout ;
wire Xd_0__inst_mult_26_24 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_10_23_sumout ;
wire Xd_0__inst_mult_10_24 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_21_23_sumout ;
wire Xd_0__inst_mult_21_24 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_14_23_sumout ;
wire Xd_0__inst_mult_14_24 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_25_23_sumout ;
wire Xd_0__inst_mult_25_24 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_87_cout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_28_23_sumout ;
wire Xd_0__inst_mult_28_24 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_30_23_sumout ;
wire Xd_0__inst_mult_30_24 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_23_23_sumout ;
wire Xd_0__inst_mult_23_24 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_2_23_sumout ;
wire Xd_0__inst_mult_2_24 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_4_23_sumout ;
wire Xd_0__inst_mult_4_24 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_6_23_sumout ;
wire Xd_0__inst_mult_6_24 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_8_23_sumout ;
wire Xd_0__inst_mult_8_24 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_9_23_sumout ;
wire Xd_0__inst_mult_9_24 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_27_23_sumout ;
wire Xd_0__inst_mult_27_24 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_29_23_sumout ;
wire Xd_0__inst_mult_29_24 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_10_28_sumout ;
wire Xd_0__inst_mult_10_29 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_31_23_sumout ;
wire Xd_0__inst_mult_31_24 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_3_23_sumout ;
wire Xd_0__inst_mult_3_24 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_5_23_sumout ;
wire Xd_0__inst_mult_5_24 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_7_23_sumout ;
wire Xd_0__inst_mult_7_24 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_82 ;
wire Xd_0__inst_mult_1_23_sumout ;
wire Xd_0__inst_mult_1_24 ;
wire Xd_0__inst_mult_5_84 ;
wire Xd_0__inst_mult_5_85 ;
wire Xd_0__inst_mult_6_84 ;
wire Xd_0__inst_mult_6_85 ;
wire Xd_0__inst_i21_1_sumout ;
wire Xd_0__inst_i21_2 ;
wire Xd_0__inst_mult_7_84 ;
wire Xd_0__inst_mult_7_85 ;
wire Xd_0__inst_mult_8_84 ;
wire Xd_0__inst_mult_8_85 ;
wire Xd_0__inst_i21_6_sumout ;
wire Xd_0__inst_i21_7 ;
wire Xd_0__inst_mult_9_84 ;
wire Xd_0__inst_mult_9_85 ;
wire Xd_0__inst_mult_20_84 ;
wire Xd_0__inst_mult_20_85 ;
wire Xd_0__inst_i21_11_sumout ;
wire Xd_0__inst_i21_12 ;
wire Xd_0__inst_mult_19_84 ;
wire Xd_0__inst_mult_19_85 ;
wire Xd_0__inst_mult_11_84 ;
wire Xd_0__inst_mult_11_85 ;
wire Xd_0__inst_i21_16_sumout ;
wire Xd_0__inst_i21_17 ;
wire Xd_0__inst_mult_18_84 ;
wire Xd_0__inst_mult_18_85 ;
wire Xd_0__inst_mult_17_84 ;
wire Xd_0__inst_mult_17_85 ;
wire Xd_0__inst_i21_21_sumout ;
wire Xd_0__inst_i21_22 ;
wire Xd_0__inst_mult_16_84 ;
wire Xd_0__inst_mult_16_85 ;
wire Xd_0__inst_mult_10_84 ;
wire Xd_0__inst_mult_10_85 ;
wire Xd_0__inst_i21_26_sumout ;
wire Xd_0__inst_i21_27 ;
wire Xd_0__inst_mult_15_84 ;
wire Xd_0__inst_mult_15_85 ;
wire Xd_0__inst_mult_14_84 ;
wire Xd_0__inst_mult_14_85 ;
wire Xd_0__inst_i21_31_sumout ;
wire Xd_0__inst_i21_32 ;
wire Xd_0__inst_mult_13_84 ;
wire Xd_0__inst_mult_13_85 ;
wire Xd_0__inst_mult_12_84 ;
wire Xd_0__inst_mult_12_85 ;
wire Xd_0__inst_i21_36_sumout ;
wire Xd_0__inst_i21_37 ;
wire Xd_0__inst_mult_31_85 ;
wire Xd_0__inst_mult_31_86 ;
wire Xd_0__inst_mult_30_85 ;
wire Xd_0__inst_mult_30_86 ;
wire Xd_0__inst_mult_29_85 ;
wire Xd_0__inst_mult_29_86 ;
wire Xd_0__inst_mult_28_85 ;
wire Xd_0__inst_mult_28_86 ;
wire Xd_0__inst_mult_27_85 ;
wire Xd_0__inst_mult_27_86 ;
wire Xd_0__inst_mult_26_85 ;
wire Xd_0__inst_mult_26_86 ;
wire Xd_0__inst_mult_25_85 ;
wire Xd_0__inst_mult_25_86 ;
wire Xd_0__inst_mult_24_85 ;
wire Xd_0__inst_mult_24_86 ;
wire Xd_0__inst_mult_23_85 ;
wire Xd_0__inst_mult_23_86 ;
wire Xd_0__inst_mult_22_85 ;
wire Xd_0__inst_mult_22_86 ;
wire Xd_0__inst_mult_21_85 ;
wire Xd_0__inst_mult_21_86 ;
wire Xd_0__inst_mult_20_89 ;
wire Xd_0__inst_mult_20_90 ;
wire Xd_0__inst_mult_19_89 ;
wire Xd_0__inst_mult_19_90 ;
wire Xd_0__inst_mult_18_89 ;
wire Xd_0__inst_mult_18_90 ;
wire Xd_0__inst_mult_17_89 ;
wire Xd_0__inst_mult_17_90 ;
wire Xd_0__inst_mult_16_89 ;
wire Xd_0__inst_mult_16_90 ;
wire Xd_0__inst_mult_15_89 ;
wire Xd_0__inst_mult_15_90 ;
wire Xd_0__inst_mult_14_89 ;
wire Xd_0__inst_mult_14_90 ;
wire Xd_0__inst_mult_13_89 ;
wire Xd_0__inst_mult_13_90 ;
wire Xd_0__inst_mult_12_89 ;
wire Xd_0__inst_mult_12_90 ;
wire Xd_0__inst_mult_11_89 ;
wire Xd_0__inst_mult_11_90 ;
wire Xd_0__inst_mult_10_89 ;
wire Xd_0__inst_mult_10_90 ;
wire Xd_0__inst_mult_9_89 ;
wire Xd_0__inst_mult_9_90 ;
wire Xd_0__inst_mult_8_89 ;
wire Xd_0__inst_mult_8_90 ;
wire Xd_0__inst_mult_7_89 ;
wire Xd_0__inst_mult_7_90 ;
wire Xd_0__inst_mult_6_89 ;
wire Xd_0__inst_mult_6_90 ;
wire Xd_0__inst_mult_5_89 ;
wire Xd_0__inst_mult_5_90 ;
wire Xd_0__inst_mult_4_85 ;
wire Xd_0__inst_mult_4_86 ;
wire Xd_0__inst_mult_3_85 ;
wire Xd_0__inst_mult_3_86 ;
wire Xd_0__inst_mult_2_85 ;
wire Xd_0__inst_mult_2_86 ;
wire Xd_0__inst_mult_1_85 ;
wire Xd_0__inst_mult_1_86 ;
wire Xd_0__inst_mult_0_85 ;
wire Xd_0__inst_mult_0_86 ;
wire Xd_0__inst_mult_31_90 ;
wire Xd_0__inst_mult_31_91 ;
wire Xd_0__inst_mult_30_90 ;
wire Xd_0__inst_mult_30_91 ;
wire Xd_0__inst_mult_29_90 ;
wire Xd_0__inst_mult_29_91 ;
wire Xd_0__inst_mult_28_90 ;
wire Xd_0__inst_mult_28_91 ;
wire Xd_0__inst_mult_27_90 ;
wire Xd_0__inst_mult_27_91 ;
wire Xd_0__inst_mult_26_90 ;
wire Xd_0__inst_mult_26_91 ;
wire Xd_0__inst_mult_25_90 ;
wire Xd_0__inst_mult_25_91 ;
wire Xd_0__inst_mult_24_90 ;
wire Xd_0__inst_mult_24_91 ;
wire Xd_0__inst_mult_23_90 ;
wire Xd_0__inst_mult_23_91 ;
wire Xd_0__inst_mult_22_90 ;
wire Xd_0__inst_mult_22_91 ;
wire Xd_0__inst_mult_21_90 ;
wire Xd_0__inst_mult_21_91 ;
wire Xd_0__inst_mult_20_93 ;
wire Xd_0__inst_mult_20_94 ;
wire Xd_0__inst_mult_19_93 ;
wire Xd_0__inst_mult_19_94 ;
wire Xd_0__inst_mult_18_93 ;
wire Xd_0__inst_mult_18_94 ;
wire Xd_0__inst_mult_17_93 ;
wire Xd_0__inst_mult_17_94 ;
wire Xd_0__inst_mult_16_93 ;
wire Xd_0__inst_mult_16_94 ;
wire Xd_0__inst_mult_15_93 ;
wire Xd_0__inst_mult_15_94 ;
wire Xd_0__inst_mult_14_93 ;
wire Xd_0__inst_mult_14_94 ;
wire Xd_0__inst_mult_13_93 ;
wire Xd_0__inst_mult_13_94 ;
wire Xd_0__inst_mult_12_93 ;
wire Xd_0__inst_mult_12_94 ;
wire Xd_0__inst_mult_11_93 ;
wire Xd_0__inst_mult_11_94 ;
wire Xd_0__inst_mult_10_93 ;
wire Xd_0__inst_mult_10_94 ;
wire Xd_0__inst_mult_9_93 ;
wire Xd_0__inst_mult_9_94 ;
wire Xd_0__inst_mult_8_93 ;
wire Xd_0__inst_mult_8_94 ;
wire Xd_0__inst_mult_7_93 ;
wire Xd_0__inst_mult_7_94 ;
wire Xd_0__inst_mult_6_93 ;
wire Xd_0__inst_mult_6_94 ;
wire Xd_0__inst_mult_5_93 ;
wire Xd_0__inst_mult_5_94 ;
wire Xd_0__inst_mult_4_90 ;
wire Xd_0__inst_mult_4_91 ;
wire Xd_0__inst_mult_3_90 ;
wire Xd_0__inst_mult_3_91 ;
wire Xd_0__inst_mult_2_90 ;
wire Xd_0__inst_mult_2_91 ;
wire Xd_0__inst_mult_1_90 ;
wire Xd_0__inst_mult_1_91 ;
wire Xd_0__inst_mult_0_90 ;
wire Xd_0__inst_mult_0_91 ;
wire Xd_0__inst_mult_31_94 ;
wire Xd_0__inst_mult_31_95 ;
wire Xd_0__inst_mult_30_94 ;
wire Xd_0__inst_mult_30_95 ;
wire Xd_0__inst_mult_29_94 ;
wire Xd_0__inst_mult_29_95 ;
wire Xd_0__inst_mult_28_94 ;
wire Xd_0__inst_mult_28_95 ;
wire Xd_0__inst_mult_27_94 ;
wire Xd_0__inst_mult_27_95 ;
wire Xd_0__inst_mult_26_94 ;
wire Xd_0__inst_mult_26_95 ;
wire Xd_0__inst_mult_25_94 ;
wire Xd_0__inst_mult_25_95 ;
wire Xd_0__inst_mult_24_94 ;
wire Xd_0__inst_mult_24_95 ;
wire Xd_0__inst_mult_23_94 ;
wire Xd_0__inst_mult_23_95 ;
wire Xd_0__inst_mult_22_94 ;
wire Xd_0__inst_mult_22_95 ;
wire Xd_0__inst_mult_21_94 ;
wire Xd_0__inst_mult_21_95 ;
wire Xd_0__inst_mult_20_98 ;
wire Xd_0__inst_mult_20_99 ;
wire Xd_0__inst_mult_19_98 ;
wire Xd_0__inst_mult_19_99 ;
wire Xd_0__inst_mult_18_98 ;
wire Xd_0__inst_mult_18_99 ;
wire Xd_0__inst_mult_17_98 ;
wire Xd_0__inst_mult_17_99 ;
wire Xd_0__inst_mult_16_98 ;
wire Xd_0__inst_mult_16_99 ;
wire Xd_0__inst_mult_15_98 ;
wire Xd_0__inst_mult_15_99 ;
wire Xd_0__inst_mult_14_98 ;
wire Xd_0__inst_mult_14_99 ;
wire Xd_0__inst_mult_13_98 ;
wire Xd_0__inst_mult_13_99 ;
wire Xd_0__inst_mult_12_98 ;
wire Xd_0__inst_mult_12_99 ;
wire Xd_0__inst_mult_11_98 ;
wire Xd_0__inst_mult_11_99 ;
wire Xd_0__inst_mult_10_98 ;
wire Xd_0__inst_mult_10_99 ;
wire Xd_0__inst_mult_9_98 ;
wire Xd_0__inst_mult_9_99 ;
wire Xd_0__inst_mult_8_98 ;
wire Xd_0__inst_mult_8_99 ;
wire Xd_0__inst_mult_7_98 ;
wire Xd_0__inst_mult_7_99 ;
wire Xd_0__inst_mult_6_98 ;
wire Xd_0__inst_mult_6_99 ;
wire Xd_0__inst_mult_5_98 ;
wire Xd_0__inst_mult_5_99 ;
wire Xd_0__inst_mult_4_94 ;
wire Xd_0__inst_mult_4_95 ;
wire Xd_0__inst_mult_3_94 ;
wire Xd_0__inst_mult_3_95 ;
wire Xd_0__inst_mult_2_94 ;
wire Xd_0__inst_mult_2_95 ;
wire Xd_0__inst_mult_1_94 ;
wire Xd_0__inst_mult_1_95 ;
wire Xd_0__inst_mult_0_94 ;
wire Xd_0__inst_mult_0_95 ;
wire Xd_0__inst_mult_31_99 ;
wire Xd_0__inst_mult_31_100 ;
wire Xd_0__inst_mult_30_99 ;
wire Xd_0__inst_mult_30_100 ;
wire Xd_0__inst_mult_29_99 ;
wire Xd_0__inst_mult_29_100 ;
wire Xd_0__inst_mult_28_99 ;
wire Xd_0__inst_mult_28_100 ;
wire Xd_0__inst_mult_27_99 ;
wire Xd_0__inst_mult_27_100 ;
wire Xd_0__inst_mult_26_99 ;
wire Xd_0__inst_mult_26_100 ;
wire Xd_0__inst_mult_25_99 ;
wire Xd_0__inst_mult_25_100 ;
wire Xd_0__inst_mult_24_99 ;
wire Xd_0__inst_mult_24_100 ;
wire Xd_0__inst_mult_23_99 ;
wire Xd_0__inst_mult_23_100 ;
wire Xd_0__inst_mult_22_99 ;
wire Xd_0__inst_mult_22_100 ;
wire Xd_0__inst_mult_21_99 ;
wire Xd_0__inst_mult_21_100 ;
wire Xd_0__inst_mult_20_103 ;
wire Xd_0__inst_mult_20_104 ;
wire Xd_0__inst_mult_19_103 ;
wire Xd_0__inst_mult_19_104 ;
wire Xd_0__inst_mult_18_103 ;
wire Xd_0__inst_mult_18_104 ;
wire Xd_0__inst_mult_17_103 ;
wire Xd_0__inst_mult_17_104 ;
wire Xd_0__inst_mult_16_103 ;
wire Xd_0__inst_mult_16_104 ;
wire Xd_0__inst_mult_15_103 ;
wire Xd_0__inst_mult_15_104 ;
wire Xd_0__inst_mult_14_103 ;
wire Xd_0__inst_mult_14_104 ;
wire Xd_0__inst_mult_13_103 ;
wire Xd_0__inst_mult_13_104 ;
wire Xd_0__inst_mult_12_103 ;
wire Xd_0__inst_mult_12_104 ;
wire Xd_0__inst_mult_11_103 ;
wire Xd_0__inst_mult_11_104 ;
wire Xd_0__inst_mult_10_103 ;
wire Xd_0__inst_mult_10_104 ;
wire Xd_0__inst_mult_9_103 ;
wire Xd_0__inst_mult_9_104 ;
wire Xd_0__inst_mult_8_103 ;
wire Xd_0__inst_mult_8_104 ;
wire Xd_0__inst_mult_7_103 ;
wire Xd_0__inst_mult_7_104 ;
wire Xd_0__inst_mult_6_103 ;
wire Xd_0__inst_mult_6_104 ;
wire Xd_0__inst_mult_5_103 ;
wire Xd_0__inst_mult_5_104 ;
wire Xd_0__inst_mult_4_99 ;
wire Xd_0__inst_mult_4_100 ;
wire Xd_0__inst_mult_3_99 ;
wire Xd_0__inst_mult_3_100 ;
wire Xd_0__inst_mult_2_99 ;
wire Xd_0__inst_mult_2_100 ;
wire Xd_0__inst_mult_1_99 ;
wire Xd_0__inst_mult_1_100 ;
wire Xd_0__inst_mult_0_99 ;
wire Xd_0__inst_mult_0_100 ;
wire Xd_0__inst_mult_31_104 ;
wire Xd_0__inst_mult_31_105 ;
wire Xd_0__inst_mult_30_104 ;
wire Xd_0__inst_mult_30_105 ;
wire Xd_0__inst_mult_29_104 ;
wire Xd_0__inst_mult_29_105 ;
wire Xd_0__inst_mult_28_104 ;
wire Xd_0__inst_mult_28_105 ;
wire Xd_0__inst_mult_27_104 ;
wire Xd_0__inst_mult_27_105 ;
wire Xd_0__inst_mult_26_104 ;
wire Xd_0__inst_mult_26_105 ;
wire Xd_0__inst_mult_25_104 ;
wire Xd_0__inst_mult_25_105 ;
wire Xd_0__inst_mult_24_104 ;
wire Xd_0__inst_mult_24_105 ;
wire Xd_0__inst_mult_23_104 ;
wire Xd_0__inst_mult_23_105 ;
wire Xd_0__inst_mult_22_104 ;
wire Xd_0__inst_mult_22_105 ;
wire Xd_0__inst_mult_21_104 ;
wire Xd_0__inst_mult_21_105 ;
wire Xd_0__inst_mult_20_108 ;
wire Xd_0__inst_mult_20_109 ;
wire Xd_0__inst_mult_19_108 ;
wire Xd_0__inst_mult_19_109 ;
wire Xd_0__inst_mult_18_108 ;
wire Xd_0__inst_mult_18_109 ;
wire Xd_0__inst_mult_17_108 ;
wire Xd_0__inst_mult_17_109 ;
wire Xd_0__inst_mult_16_108 ;
wire Xd_0__inst_mult_16_109 ;
wire Xd_0__inst_mult_15_108 ;
wire Xd_0__inst_mult_15_109 ;
wire Xd_0__inst_mult_14_108 ;
wire Xd_0__inst_mult_14_109 ;
wire Xd_0__inst_mult_13_108 ;
wire Xd_0__inst_mult_13_109 ;
wire Xd_0__inst_mult_12_108 ;
wire Xd_0__inst_mult_12_109 ;
wire Xd_0__inst_mult_11_108 ;
wire Xd_0__inst_mult_11_109 ;
wire Xd_0__inst_mult_10_108 ;
wire Xd_0__inst_mult_10_109 ;
wire Xd_0__inst_mult_9_108 ;
wire Xd_0__inst_mult_9_109 ;
wire Xd_0__inst_mult_8_108 ;
wire Xd_0__inst_mult_8_109 ;
wire Xd_0__inst_mult_7_108 ;
wire Xd_0__inst_mult_7_109 ;
wire Xd_0__inst_mult_6_108 ;
wire Xd_0__inst_mult_6_109 ;
wire Xd_0__inst_mult_5_108 ;
wire Xd_0__inst_mult_5_109 ;
wire Xd_0__inst_mult_4_104 ;
wire Xd_0__inst_mult_4_105 ;
wire Xd_0__inst_mult_3_104 ;
wire Xd_0__inst_mult_3_105 ;
wire Xd_0__inst_mult_2_104 ;
wire Xd_0__inst_mult_2_105 ;
wire Xd_0__inst_mult_1_104 ;
wire Xd_0__inst_mult_1_105 ;
wire Xd_0__inst_mult_0_104 ;
wire Xd_0__inst_mult_0_105 ;
wire Xd_0__inst_mult_31_109 ;
wire Xd_0__inst_mult_31_110 ;
wire Xd_0__inst_mult_30_109 ;
wire Xd_0__inst_mult_30_110 ;
wire Xd_0__inst_mult_29_109 ;
wire Xd_0__inst_mult_29_110 ;
wire Xd_0__inst_mult_28_109 ;
wire Xd_0__inst_mult_28_110 ;
wire Xd_0__inst_mult_27_109 ;
wire Xd_0__inst_mult_27_110 ;
wire Xd_0__inst_mult_26_109 ;
wire Xd_0__inst_mult_26_110 ;
wire Xd_0__inst_mult_25_109 ;
wire Xd_0__inst_mult_25_110 ;
wire Xd_0__inst_mult_24_109 ;
wire Xd_0__inst_mult_24_110 ;
wire Xd_0__inst_mult_23_109 ;
wire Xd_0__inst_mult_23_110 ;
wire Xd_0__inst_mult_22_109 ;
wire Xd_0__inst_mult_22_110 ;
wire Xd_0__inst_mult_21_109 ;
wire Xd_0__inst_mult_21_110 ;
wire Xd_0__inst_mult_20_113 ;
wire Xd_0__inst_mult_20_114 ;
wire Xd_0__inst_mult_19_113 ;
wire Xd_0__inst_mult_19_114 ;
wire Xd_0__inst_mult_18_113 ;
wire Xd_0__inst_mult_18_114 ;
wire Xd_0__inst_mult_17_113 ;
wire Xd_0__inst_mult_17_114 ;
wire Xd_0__inst_mult_16_113 ;
wire Xd_0__inst_mult_16_114 ;
wire Xd_0__inst_mult_15_113 ;
wire Xd_0__inst_mult_15_114 ;
wire Xd_0__inst_mult_14_113 ;
wire Xd_0__inst_mult_14_114 ;
wire Xd_0__inst_mult_13_113 ;
wire Xd_0__inst_mult_13_114 ;
wire Xd_0__inst_mult_12_113 ;
wire Xd_0__inst_mult_12_114 ;
wire Xd_0__inst_mult_11_113 ;
wire Xd_0__inst_mult_11_114 ;
wire Xd_0__inst_mult_10_113 ;
wire Xd_0__inst_mult_10_114 ;
wire Xd_0__inst_mult_9_113 ;
wire Xd_0__inst_mult_9_114 ;
wire Xd_0__inst_mult_8_113 ;
wire Xd_0__inst_mult_8_114 ;
wire Xd_0__inst_mult_7_113 ;
wire Xd_0__inst_mult_7_114 ;
wire Xd_0__inst_mult_6_113 ;
wire Xd_0__inst_mult_6_114 ;
wire Xd_0__inst_mult_5_113 ;
wire Xd_0__inst_mult_5_114 ;
wire Xd_0__inst_mult_4_109 ;
wire Xd_0__inst_mult_4_110 ;
wire Xd_0__inst_mult_3_109 ;
wire Xd_0__inst_mult_3_110 ;
wire Xd_0__inst_mult_2_109 ;
wire Xd_0__inst_mult_2_110 ;
wire Xd_0__inst_mult_1_109 ;
wire Xd_0__inst_mult_1_110 ;
wire Xd_0__inst_mult_0_109 ;
wire Xd_0__inst_mult_0_110 ;
wire Xd_0__inst_mult_31_114 ;
wire Xd_0__inst_mult_31_115 ;
wire Xd_0__inst_mult_30_114 ;
wire Xd_0__inst_mult_30_115 ;
wire Xd_0__inst_mult_29_114 ;
wire Xd_0__inst_mult_29_115 ;
wire Xd_0__inst_mult_28_114 ;
wire Xd_0__inst_mult_28_115 ;
wire Xd_0__inst_mult_27_114 ;
wire Xd_0__inst_mult_27_115 ;
wire Xd_0__inst_mult_26_114 ;
wire Xd_0__inst_mult_26_115 ;
wire Xd_0__inst_mult_25_114 ;
wire Xd_0__inst_mult_25_115 ;
wire Xd_0__inst_mult_24_114 ;
wire Xd_0__inst_mult_24_115 ;
wire Xd_0__inst_mult_23_114 ;
wire Xd_0__inst_mult_23_115 ;
wire Xd_0__inst_mult_22_114 ;
wire Xd_0__inst_mult_22_115 ;
wire Xd_0__inst_mult_21_114 ;
wire Xd_0__inst_mult_21_115 ;
wire Xd_0__inst_mult_20_118 ;
wire Xd_0__inst_mult_20_119 ;
wire Xd_0__inst_mult_19_118 ;
wire Xd_0__inst_mult_19_119 ;
wire Xd_0__inst_mult_18_118 ;
wire Xd_0__inst_mult_18_119 ;
wire Xd_0__inst_mult_17_118 ;
wire Xd_0__inst_mult_17_119 ;
wire Xd_0__inst_mult_16_118 ;
wire Xd_0__inst_mult_16_119 ;
wire Xd_0__inst_mult_15_118 ;
wire Xd_0__inst_mult_15_119 ;
wire Xd_0__inst_mult_14_118 ;
wire Xd_0__inst_mult_14_119 ;
wire Xd_0__inst_mult_13_118 ;
wire Xd_0__inst_mult_13_119 ;
wire Xd_0__inst_mult_12_118 ;
wire Xd_0__inst_mult_12_119 ;
wire Xd_0__inst_mult_11_118 ;
wire Xd_0__inst_mult_11_119 ;
wire Xd_0__inst_mult_10_118 ;
wire Xd_0__inst_mult_10_119 ;
wire Xd_0__inst_mult_9_118 ;
wire Xd_0__inst_mult_9_119 ;
wire Xd_0__inst_mult_8_118 ;
wire Xd_0__inst_mult_8_119 ;
wire Xd_0__inst_mult_7_118 ;
wire Xd_0__inst_mult_7_119 ;
wire Xd_0__inst_mult_6_118 ;
wire Xd_0__inst_mult_6_119 ;
wire Xd_0__inst_mult_5_118 ;
wire Xd_0__inst_mult_5_119 ;
wire Xd_0__inst_mult_4_114 ;
wire Xd_0__inst_mult_4_115 ;
wire Xd_0__inst_mult_3_114 ;
wire Xd_0__inst_mult_3_115 ;
wire Xd_0__inst_mult_2_114 ;
wire Xd_0__inst_mult_2_115 ;
wire Xd_0__inst_mult_1_114 ;
wire Xd_0__inst_mult_1_115 ;
wire Xd_0__inst_mult_0_114 ;
wire Xd_0__inst_mult_0_115 ;
wire Xd_0__inst_mult_31_119 ;
wire Xd_0__inst_mult_31_120 ;
wire Xd_0__inst_mult_30_119 ;
wire Xd_0__inst_mult_30_120 ;
wire Xd_0__inst_mult_29_119 ;
wire Xd_0__inst_mult_29_120 ;
wire Xd_0__inst_mult_28_119 ;
wire Xd_0__inst_mult_28_120 ;
wire Xd_0__inst_mult_27_119 ;
wire Xd_0__inst_mult_27_120 ;
wire Xd_0__inst_mult_26_119 ;
wire Xd_0__inst_mult_26_120 ;
wire Xd_0__inst_mult_25_119 ;
wire Xd_0__inst_mult_25_120 ;
wire Xd_0__inst_mult_24_119 ;
wire Xd_0__inst_mult_24_120 ;
wire Xd_0__inst_mult_23_119 ;
wire Xd_0__inst_mult_23_120 ;
wire Xd_0__inst_mult_22_119 ;
wire Xd_0__inst_mult_22_120 ;
wire Xd_0__inst_mult_21_119 ;
wire Xd_0__inst_mult_21_120 ;
wire Xd_0__inst_mult_20_123 ;
wire Xd_0__inst_mult_20_124 ;
wire Xd_0__inst_mult_19_123 ;
wire Xd_0__inst_mult_19_124 ;
wire Xd_0__inst_mult_18_123 ;
wire Xd_0__inst_mult_18_124 ;
wire Xd_0__inst_mult_17_123 ;
wire Xd_0__inst_mult_17_124 ;
wire Xd_0__inst_mult_16_123 ;
wire Xd_0__inst_mult_16_124 ;
wire Xd_0__inst_mult_15_123 ;
wire Xd_0__inst_mult_15_124 ;
wire Xd_0__inst_mult_14_123 ;
wire Xd_0__inst_mult_14_124 ;
wire Xd_0__inst_mult_13_123 ;
wire Xd_0__inst_mult_13_124 ;
wire Xd_0__inst_mult_12_123 ;
wire Xd_0__inst_mult_12_124 ;
wire Xd_0__inst_mult_11_123 ;
wire Xd_0__inst_mult_11_124 ;
wire Xd_0__inst_mult_10_123 ;
wire Xd_0__inst_mult_10_124 ;
wire Xd_0__inst_mult_9_123 ;
wire Xd_0__inst_mult_9_124 ;
wire Xd_0__inst_mult_8_123 ;
wire Xd_0__inst_mult_8_124 ;
wire Xd_0__inst_mult_7_123 ;
wire Xd_0__inst_mult_7_124 ;
wire Xd_0__inst_mult_6_123 ;
wire Xd_0__inst_mult_6_124 ;
wire Xd_0__inst_mult_5_123 ;
wire Xd_0__inst_mult_5_124 ;
wire Xd_0__inst_mult_4_119 ;
wire Xd_0__inst_mult_4_120 ;
wire Xd_0__inst_mult_3_119 ;
wire Xd_0__inst_mult_3_120 ;
wire Xd_0__inst_mult_2_119 ;
wire Xd_0__inst_mult_2_120 ;
wire Xd_0__inst_mult_1_119 ;
wire Xd_0__inst_mult_1_120 ;
wire Xd_0__inst_mult_0_119 ;
wire Xd_0__inst_mult_0_120 ;
wire Xd_0__inst_mult_31_124 ;
wire Xd_0__inst_mult_31_125 ;
wire Xd_0__inst_mult_30_124 ;
wire Xd_0__inst_mult_30_125 ;
wire Xd_0__inst_mult_29_124 ;
wire Xd_0__inst_mult_29_125 ;
wire Xd_0__inst_mult_28_124 ;
wire Xd_0__inst_mult_28_125 ;
wire Xd_0__inst_mult_27_124 ;
wire Xd_0__inst_mult_27_125 ;
wire Xd_0__inst_mult_26_124 ;
wire Xd_0__inst_mult_26_125 ;
wire Xd_0__inst_mult_25_124 ;
wire Xd_0__inst_mult_25_125 ;
wire Xd_0__inst_mult_24_124 ;
wire Xd_0__inst_mult_24_125 ;
wire Xd_0__inst_mult_23_124 ;
wire Xd_0__inst_mult_23_125 ;
wire Xd_0__inst_mult_22_124 ;
wire Xd_0__inst_mult_22_125 ;
wire Xd_0__inst_mult_21_124 ;
wire Xd_0__inst_mult_21_125 ;
wire Xd_0__inst_mult_20_128 ;
wire Xd_0__inst_mult_20_129 ;
wire Xd_0__inst_mult_19_128 ;
wire Xd_0__inst_mult_19_129 ;
wire Xd_0__inst_mult_18_128 ;
wire Xd_0__inst_mult_18_129 ;
wire Xd_0__inst_mult_17_128 ;
wire Xd_0__inst_mult_17_129 ;
wire Xd_0__inst_mult_16_128 ;
wire Xd_0__inst_mult_16_129 ;
wire Xd_0__inst_mult_15_128 ;
wire Xd_0__inst_mult_15_129 ;
wire Xd_0__inst_mult_14_128 ;
wire Xd_0__inst_mult_14_129 ;
wire Xd_0__inst_mult_13_128 ;
wire Xd_0__inst_mult_13_129 ;
wire Xd_0__inst_mult_12_128 ;
wire Xd_0__inst_mult_12_129 ;
wire Xd_0__inst_mult_11_128 ;
wire Xd_0__inst_mult_11_129 ;
wire Xd_0__inst_mult_10_128 ;
wire Xd_0__inst_mult_10_129 ;
wire Xd_0__inst_mult_9_128 ;
wire Xd_0__inst_mult_9_129 ;
wire Xd_0__inst_mult_8_128 ;
wire Xd_0__inst_mult_8_129 ;
wire Xd_0__inst_mult_7_128 ;
wire Xd_0__inst_mult_7_129 ;
wire Xd_0__inst_mult_6_128 ;
wire Xd_0__inst_mult_6_129 ;
wire Xd_0__inst_mult_5_128 ;
wire Xd_0__inst_mult_5_129 ;
wire Xd_0__inst_mult_4_124 ;
wire Xd_0__inst_mult_4_125 ;
wire Xd_0__inst_mult_3_124 ;
wire Xd_0__inst_mult_3_125 ;
wire Xd_0__inst_mult_2_124 ;
wire Xd_0__inst_mult_2_125 ;
wire Xd_0__inst_mult_1_124 ;
wire Xd_0__inst_mult_1_125 ;
wire Xd_0__inst_mult_0_124 ;
wire Xd_0__inst_mult_0_125 ;
wire Xd_0__inst_mult_31_129 ;
wire Xd_0__inst_mult_31_130 ;
wire Xd_0__inst_mult_30_129 ;
wire Xd_0__inst_mult_30_130 ;
wire Xd_0__inst_mult_29_129 ;
wire Xd_0__inst_mult_29_130 ;
wire Xd_0__inst_mult_28_129 ;
wire Xd_0__inst_mult_28_130 ;
wire Xd_0__inst_mult_27_129 ;
wire Xd_0__inst_mult_27_130 ;
wire Xd_0__inst_mult_26_129 ;
wire Xd_0__inst_mult_26_130 ;
wire Xd_0__inst_mult_25_129 ;
wire Xd_0__inst_mult_25_130 ;
wire Xd_0__inst_mult_24_129 ;
wire Xd_0__inst_mult_24_130 ;
wire Xd_0__inst_mult_23_129 ;
wire Xd_0__inst_mult_23_130 ;
wire Xd_0__inst_mult_22_129 ;
wire Xd_0__inst_mult_22_130 ;
wire Xd_0__inst_mult_21_129 ;
wire Xd_0__inst_mult_21_130 ;
wire Xd_0__inst_mult_20_133 ;
wire Xd_0__inst_mult_20_134 ;
wire Xd_0__inst_mult_19_133 ;
wire Xd_0__inst_mult_19_134 ;
wire Xd_0__inst_mult_18_133 ;
wire Xd_0__inst_mult_18_134 ;
wire Xd_0__inst_mult_17_133 ;
wire Xd_0__inst_mult_17_134 ;
wire Xd_0__inst_mult_16_133 ;
wire Xd_0__inst_mult_16_134 ;
wire Xd_0__inst_mult_15_133 ;
wire Xd_0__inst_mult_15_134 ;
wire Xd_0__inst_mult_14_133 ;
wire Xd_0__inst_mult_14_134 ;
wire Xd_0__inst_mult_13_133 ;
wire Xd_0__inst_mult_13_134 ;
wire Xd_0__inst_mult_12_133 ;
wire Xd_0__inst_mult_12_134 ;
wire Xd_0__inst_mult_11_133 ;
wire Xd_0__inst_mult_11_134 ;
wire Xd_0__inst_mult_10_133 ;
wire Xd_0__inst_mult_10_134 ;
wire Xd_0__inst_mult_9_133 ;
wire Xd_0__inst_mult_9_134 ;
wire Xd_0__inst_mult_8_133 ;
wire Xd_0__inst_mult_8_134 ;
wire Xd_0__inst_mult_7_133 ;
wire Xd_0__inst_mult_7_134 ;
wire Xd_0__inst_mult_6_133 ;
wire Xd_0__inst_mult_6_134 ;
wire Xd_0__inst_mult_5_133 ;
wire Xd_0__inst_mult_5_134 ;
wire Xd_0__inst_mult_4_129 ;
wire Xd_0__inst_mult_4_130 ;
wire Xd_0__inst_mult_3_129 ;
wire Xd_0__inst_mult_3_130 ;
wire Xd_0__inst_mult_2_129 ;
wire Xd_0__inst_mult_2_130 ;
wire Xd_0__inst_mult_1_129 ;
wire Xd_0__inst_mult_1_130 ;
wire Xd_0__inst_mult_0_129 ;
wire Xd_0__inst_mult_0_130 ;
wire Xd_0__inst_mult_31_134 ;
wire Xd_0__inst_mult_30_134 ;
wire Xd_0__inst_mult_29_134 ;
wire Xd_0__inst_mult_28_134 ;
wire Xd_0__inst_mult_27_134 ;
wire Xd_0__inst_mult_26_134 ;
wire Xd_0__inst_mult_25_134 ;
wire Xd_0__inst_mult_24_134 ;
wire Xd_0__inst_mult_23_134 ;
wire Xd_0__inst_mult_22_134 ;
wire Xd_0__inst_mult_21_134 ;
wire Xd_0__inst_mult_20_138 ;
wire Xd_0__inst_mult_19_138 ;
wire Xd_0__inst_mult_18_138 ;
wire Xd_0__inst_mult_17_138 ;
wire Xd_0__inst_mult_16_138 ;
wire Xd_0__inst_mult_15_138 ;
wire Xd_0__inst_mult_14_138 ;
wire Xd_0__inst_mult_13_138 ;
wire Xd_0__inst_mult_12_138 ;
wire Xd_0__inst_mult_11_138 ;
wire Xd_0__inst_mult_10_138 ;
wire Xd_0__inst_mult_9_138 ;
wire Xd_0__inst_mult_8_138 ;
wire Xd_0__inst_mult_7_138 ;
wire Xd_0__inst_mult_6_138 ;
wire Xd_0__inst_mult_5_138 ;
wire Xd_0__inst_mult_4_134 ;
wire Xd_0__inst_mult_3_134 ;
wire Xd_0__inst_mult_2_134 ;
wire Xd_0__inst_mult_1_134 ;
wire Xd_0__inst_mult_0_134 ;
wire Xd_0__inst_i21_41_sumout ;
wire Xd_0__inst_i21_42 ;
wire Xd_0__inst_mult_31_139 ;
wire Xd_0__inst_mult_31_140 ;
wire Xd_0__inst_mult_30_139 ;
wire Xd_0__inst_mult_30_140 ;
wire Xd_0__inst_mult_5_143 ;
wire Xd_0__inst_mult_5_144 ;
wire Xd_0__inst_i21_46_sumout ;
wire Xd_0__inst_i21_47 ;
wire Xd_0__inst_i21_51_sumout ;
wire Xd_0__inst_i21_52 ;
wire Xd_0__inst_mult_29_139 ;
wire Xd_0__inst_mult_29_140 ;
wire Xd_0__inst_mult_28_139 ;
wire Xd_0__inst_mult_28_140 ;
wire Xd_0__inst_mult_6_143 ;
wire Xd_0__inst_mult_6_144 ;
wire Xd_0__inst_i21_56_sumout ;
wire Xd_0__inst_i21_57 ;
wire Xd_0__inst_i21_61_sumout ;
wire Xd_0__inst_i21_62 ;
wire Xd_0__inst_mult_27_139 ;
wire Xd_0__inst_mult_27_140 ;
wire Xd_0__inst_mult_26_139 ;
wire Xd_0__inst_mult_26_140 ;
wire Xd_0__inst_mult_7_143 ;
wire Xd_0__inst_mult_7_144 ;
wire Xd_0__inst_i21_66_sumout ;
wire Xd_0__inst_i21_67 ;
wire Xd_0__inst_i21_71_sumout ;
wire Xd_0__inst_i21_72 ;
wire Xd_0__inst_mult_25_139 ;
wire Xd_0__inst_mult_25_140 ;
wire Xd_0__inst_mult_24_139 ;
wire Xd_0__inst_mult_24_140 ;
wire Xd_0__inst_mult_8_143 ;
wire Xd_0__inst_mult_8_144 ;
wire Xd_0__inst_i21_76_sumout ;
wire Xd_0__inst_i21_77 ;
wire Xd_0__inst_mult_23_139 ;
wire Xd_0__inst_mult_23_140 ;
wire Xd_0__inst_mult_22_139 ;
wire Xd_0__inst_mult_22_140 ;
wire Xd_0__inst_mult_9_143 ;
wire Xd_0__inst_mult_9_144 ;
wire Xd_0__inst_i21_81_sumout ;
wire Xd_0__inst_i21_82 ;
wire Xd_0__inst_i21_86_sumout ;
wire Xd_0__inst_i21_87 ;
wire Xd_0__inst_mult_21_139 ;
wire Xd_0__inst_mult_21_140 ;
wire Xd_0__inst_mult_20_143 ;
wire Xd_0__inst_mult_20_144 ;
wire Xd_0__inst_mult_20_148 ;
wire Xd_0__inst_mult_20_149 ;
wire Xd_0__inst_mult_19_143 ;
wire Xd_0__inst_mult_19_144 ;
wire Xd_0__inst_mult_18_143 ;
wire Xd_0__inst_mult_18_144 ;
wire Xd_0__inst_mult_19_148 ;
wire Xd_0__inst_mult_19_149 ;
wire Xd_0__inst_i21_91_sumout ;
wire Xd_0__inst_i21_92 ;
wire Xd_0__inst_i21_96_sumout ;
wire Xd_0__inst_i21_97 ;
wire Xd_0__inst_mult_17_143 ;
wire Xd_0__inst_mult_17_144 ;
wire Xd_0__inst_mult_16_143 ;
wire Xd_0__inst_mult_16_144 ;
wire Xd_0__inst_mult_11_143 ;
wire Xd_0__inst_mult_11_144 ;
wire Xd_0__inst_i21_101_sumout ;
wire Xd_0__inst_i21_102 ;
wire Xd_0__inst_mult_15_143 ;
wire Xd_0__inst_mult_15_144 ;
wire Xd_0__inst_mult_14_143 ;
wire Xd_0__inst_mult_14_144 ;
wire Xd_0__inst_mult_18_148 ;
wire Xd_0__inst_mult_18_149 ;
wire Xd_0__inst_i21_106_sumout ;
wire Xd_0__inst_i21_107 ;
wire Xd_0__inst_i21_111_sumout ;
wire Xd_0__inst_i21_112 ;
wire Xd_0__inst_mult_13_143 ;
wire Xd_0__inst_mult_13_144 ;
wire Xd_0__inst_mult_12_143 ;
wire Xd_0__inst_mult_12_144 ;
wire Xd_0__inst_mult_17_148 ;
wire Xd_0__inst_mult_17_149 ;
wire Xd_0__inst_i21_116_sumout ;
wire Xd_0__inst_i21_117 ;
wire Xd_0__inst_mult_11_148 ;
wire Xd_0__inst_mult_11_149 ;
wire Xd_0__inst_mult_10_143 ;
wire Xd_0__inst_mult_10_144 ;
wire Xd_0__inst_mult_16_148 ;
wire Xd_0__inst_mult_16_149 ;
wire Xd_0__inst_i21_121_sumout ;
wire Xd_0__inst_i21_122 ;
wire Xd_0__inst_i21_126_sumout ;
wire Xd_0__inst_i21_127 ;
wire Xd_0__inst_mult_9_148 ;
wire Xd_0__inst_mult_9_149 ;
wire Xd_0__inst_mult_8_148 ;
wire Xd_0__inst_mult_8_149 ;
wire Xd_0__inst_mult_10_148 ;
wire Xd_0__inst_mult_10_149 ;
wire Xd_0__inst_i21_131_sumout ;
wire Xd_0__inst_i21_132 ;
wire Xd_0__inst_mult_7_148 ;
wire Xd_0__inst_mult_7_149 ;
wire Xd_0__inst_mult_6_148 ;
wire Xd_0__inst_mult_6_149 ;
wire Xd_0__inst_mult_15_148 ;
wire Xd_0__inst_mult_15_149 ;
wire Xd_0__inst_i21_136_sumout ;
wire Xd_0__inst_i21_137 ;
wire Xd_0__inst_i21_141_sumout ;
wire Xd_0__inst_i21_142 ;
wire Xd_0__inst_mult_5_148 ;
wire Xd_0__inst_mult_5_149 ;
wire Xd_0__inst_mult_4_139 ;
wire Xd_0__inst_mult_4_140 ;
wire Xd_0__inst_mult_14_148 ;
wire Xd_0__inst_mult_14_149 ;
wire Xd_0__inst_i21_146_sumout ;
wire Xd_0__inst_i21_147 ;
wire Xd_0__inst_mult_3_139 ;
wire Xd_0__inst_mult_3_140 ;
wire Xd_0__inst_mult_2_139 ;
wire Xd_0__inst_mult_2_140 ;
wire Xd_0__inst_mult_13_148 ;
wire Xd_0__inst_mult_13_149 ;
wire Xd_0__inst_i21_151_sumout ;
wire Xd_0__inst_i21_152 ;
wire Xd_0__inst_i21_156_sumout ;
wire Xd_0__inst_i21_157 ;
wire Xd_0__inst_mult_1_139 ;
wire Xd_0__inst_mult_1_140 ;
wire Xd_0__inst_mult_0_139 ;
wire Xd_0__inst_mult_0_140 ;
wire Xd_0__inst_mult_12_148 ;
wire Xd_0__inst_mult_12_149 ;
wire Xd_0__inst_mult_31_144 ;
wire Xd_0__inst_mult_31_145 ;
wire Xd_0__inst_mult_30_144 ;
wire Xd_0__inst_mult_30_145 ;
wire Xd_0__inst_mult_29_144 ;
wire Xd_0__inst_mult_29_145 ;
wire Xd_0__inst_mult_28_144 ;
wire Xd_0__inst_mult_28_145 ;
wire Xd_0__inst_mult_27_144 ;
wire Xd_0__inst_mult_27_145 ;
wire Xd_0__inst_mult_26_144 ;
wire Xd_0__inst_mult_26_145 ;
wire Xd_0__inst_mult_25_144 ;
wire Xd_0__inst_mult_25_145 ;
wire Xd_0__inst_mult_24_144 ;
wire Xd_0__inst_mult_24_145 ;
wire Xd_0__inst_mult_23_144 ;
wire Xd_0__inst_mult_23_145 ;
wire Xd_0__inst_mult_22_144 ;
wire Xd_0__inst_mult_22_145 ;
wire Xd_0__inst_mult_21_144 ;
wire Xd_0__inst_mult_21_145 ;
wire Xd_0__inst_mult_20_153 ;
wire Xd_0__inst_mult_20_154 ;
wire Xd_0__inst_mult_19_153 ;
wire Xd_0__inst_mult_19_154 ;
wire Xd_0__inst_mult_18_153 ;
wire Xd_0__inst_mult_18_154 ;
wire Xd_0__inst_mult_17_153 ;
wire Xd_0__inst_mult_17_154 ;
wire Xd_0__inst_mult_16_153 ;
wire Xd_0__inst_mult_16_154 ;
wire Xd_0__inst_mult_15_153 ;
wire Xd_0__inst_mult_15_154 ;
wire Xd_0__inst_mult_14_153 ;
wire Xd_0__inst_mult_14_154 ;
wire Xd_0__inst_mult_13_153 ;
wire Xd_0__inst_mult_13_154 ;
wire Xd_0__inst_mult_12_153 ;
wire Xd_0__inst_mult_12_154 ;
wire Xd_0__inst_mult_11_153 ;
wire Xd_0__inst_mult_11_154 ;
wire Xd_0__inst_mult_10_153 ;
wire Xd_0__inst_mult_10_154 ;
wire Xd_0__inst_mult_9_153 ;
wire Xd_0__inst_mult_9_154 ;
wire Xd_0__inst_mult_8_153 ;
wire Xd_0__inst_mult_8_154 ;
wire Xd_0__inst_mult_7_153 ;
wire Xd_0__inst_mult_7_154 ;
wire Xd_0__inst_mult_6_153 ;
wire Xd_0__inst_mult_6_154 ;
wire Xd_0__inst_mult_5_153 ;
wire Xd_0__inst_mult_5_154 ;
wire Xd_0__inst_mult_4_144 ;
wire Xd_0__inst_mult_4_145 ;
wire Xd_0__inst_mult_3_144 ;
wire Xd_0__inst_mult_3_145 ;
wire Xd_0__inst_mult_2_144 ;
wire Xd_0__inst_mult_2_145 ;
wire Xd_0__inst_mult_1_144 ;
wire Xd_0__inst_mult_1_145 ;
wire Xd_0__inst_mult_0_144 ;
wire Xd_0__inst_mult_0_145 ;
wire Xd_0__inst_mult_31_149 ;
wire Xd_0__inst_mult_31_150 ;
wire Xd_0__inst_mult_30_149 ;
wire Xd_0__inst_mult_30_150 ;
wire Xd_0__inst_mult_29_149 ;
wire Xd_0__inst_mult_29_150 ;
wire Xd_0__inst_mult_28_149 ;
wire Xd_0__inst_mult_28_150 ;
wire Xd_0__inst_mult_27_149 ;
wire Xd_0__inst_mult_27_150 ;
wire Xd_0__inst_mult_26_149 ;
wire Xd_0__inst_mult_26_150 ;
wire Xd_0__inst_mult_25_149 ;
wire Xd_0__inst_mult_25_150 ;
wire Xd_0__inst_mult_24_149 ;
wire Xd_0__inst_mult_24_150 ;
wire Xd_0__inst_mult_23_149 ;
wire Xd_0__inst_mult_23_150 ;
wire Xd_0__inst_mult_22_149 ;
wire Xd_0__inst_mult_22_150 ;
wire Xd_0__inst_mult_21_149 ;
wire Xd_0__inst_mult_21_150 ;
wire Xd_0__inst_mult_20_158 ;
wire Xd_0__inst_mult_20_159 ;
wire Xd_0__inst_mult_19_158 ;
wire Xd_0__inst_mult_19_159 ;
wire Xd_0__inst_mult_18_158 ;
wire Xd_0__inst_mult_18_159 ;
wire Xd_0__inst_mult_17_158 ;
wire Xd_0__inst_mult_17_159 ;
wire Xd_0__inst_mult_16_158 ;
wire Xd_0__inst_mult_16_159 ;
wire Xd_0__inst_mult_15_158 ;
wire Xd_0__inst_mult_15_159 ;
wire Xd_0__inst_mult_14_158 ;
wire Xd_0__inst_mult_14_159 ;
wire Xd_0__inst_mult_13_158 ;
wire Xd_0__inst_mult_13_159 ;
wire Xd_0__inst_mult_12_158 ;
wire Xd_0__inst_mult_12_159 ;
wire Xd_0__inst_mult_11_158 ;
wire Xd_0__inst_mult_11_159 ;
wire Xd_0__inst_mult_10_158 ;
wire Xd_0__inst_mult_10_159 ;
wire Xd_0__inst_mult_9_158 ;
wire Xd_0__inst_mult_9_159 ;
wire Xd_0__inst_mult_8_158 ;
wire Xd_0__inst_mult_8_159 ;
wire Xd_0__inst_mult_7_158 ;
wire Xd_0__inst_mult_7_159 ;
wire Xd_0__inst_mult_6_158 ;
wire Xd_0__inst_mult_6_159 ;
wire Xd_0__inst_mult_5_158 ;
wire Xd_0__inst_mult_5_159 ;
wire Xd_0__inst_mult_4_149 ;
wire Xd_0__inst_mult_4_150 ;
wire Xd_0__inst_mult_3_149 ;
wire Xd_0__inst_mult_3_150 ;
wire Xd_0__inst_mult_2_149 ;
wire Xd_0__inst_mult_2_150 ;
wire Xd_0__inst_mult_1_149 ;
wire Xd_0__inst_mult_1_150 ;
wire Xd_0__inst_mult_0_149 ;
wire Xd_0__inst_mult_0_150 ;
wire Xd_0__inst_mult_23_154 ;
wire Xd_0__inst_mult_23_155 ;
wire Xd_0__inst_mult_22_154 ;
wire Xd_0__inst_mult_22_155 ;
wire Xd_0__inst_mult_21_154 ;
wire Xd_0__inst_mult_21_155 ;
wire Xd_0__inst_mult_20_163 ;
wire Xd_0__inst_mult_20_164 ;
wire Xd_0__inst_mult_25_154 ;
wire Xd_0__inst_mult_25_155 ;
wire Xd_0__inst_mult_19_163 ;
wire Xd_0__inst_mult_19_164 ;
wire Xd_0__inst_mult_18_163 ;
wire Xd_0__inst_mult_18_164 ;
wire Xd_0__inst_mult_17_163 ;
wire Xd_0__inst_mult_17_164 ;
wire Xd_0__inst_mult_24_154 ;
wire Xd_0__inst_mult_24_155 ;
wire Xd_0__inst_mult_4_154 ;
wire Xd_0__inst_mult_4_155 ;
wire Xd_0__inst_mult_26_154 ;
wire Xd_0__inst_mult_26_155 ;
wire Xd_0__inst_mult_16_163 ;
wire Xd_0__inst_mult_16_164 ;
wire Xd_0__inst_mult_12_163 ;
wire Xd_0__inst_mult_12_164 ;
wire Xd_0__inst_mult_23_159 ;
wire Xd_0__inst_mult_23_160 ;
wire Xd_0__inst_mult_5_163 ;
wire Xd_0__inst_mult_5_164 ;
wire Xd_0__inst_mult_6_163 ;
wire Xd_0__inst_mult_6_164 ;
wire Xd_0__inst_mult_7_163 ;
wire Xd_0__inst_mult_7_164 ;
wire Xd_0__inst_mult_8_163 ;
wire Xd_0__inst_mult_8_164 ;
wire Xd_0__inst_mult_9_163 ;
wire Xd_0__inst_mult_9_164 ;
wire Xd_0__inst_mult_19_168 ;
wire Xd_0__inst_mult_19_169 ;
wire Xd_0__inst_mult_10_163 ;
wire Xd_0__inst_mult_10_164 ;
wire Xd_0__inst_mult_11_163 ;
wire Xd_0__inst_mult_11_164 ;
wire Xd_0__inst_mult_13_163 ;
wire Xd_0__inst_mult_13_164 ;
wire Xd_0__inst_mult_14_163 ;
wire Xd_0__inst_mult_14_164 ;
wire Xd_0__inst_mult_15_163 ;
wire Xd_0__inst_mult_15_164 ;
wire Xd_0__inst_mult_16_168 ;
wire Xd_0__inst_mult_16_169 ;
wire Xd_0__inst_mult_17_168 ;
wire Xd_0__inst_mult_17_169 ;
wire Xd_0__inst_mult_18_168 ;
wire Xd_0__inst_mult_18_169 ;
wire Xd_0__inst_mult_30_154 ;
wire Xd_0__inst_mult_30_155 ;
wire Xd_0__inst_mult_20_168 ;
wire Xd_0__inst_mult_20_169 ;
wire Xd_0__inst_mult_21_159 ;
wire Xd_0__inst_mult_21_160 ;
wire Xd_0__inst_mult_22_159 ;
wire Xd_0__inst_mult_22_160 ;
wire Xd_0__inst_mult_5_168 ;
wire Xd_0__inst_mult_5_169 ;
wire Xd_0__inst_mult_6_168 ;
wire Xd_0__inst_mult_6_169 ;
wire Xd_0__inst_mult_7_168 ;
wire Xd_0__inst_mult_7_169 ;
wire Xd_0__inst_mult_8_168 ;
wire Xd_0__inst_mult_8_169 ;
wire Xd_0__inst_mult_9_168 ;
wire Xd_0__inst_mult_9_169 ;
wire Xd_0__inst_mult_20_173 ;
wire Xd_0__inst_mult_20_174 ;
wire Xd_0__inst_mult_19_173 ;
wire Xd_0__inst_mult_19_174 ;
wire Xd_0__inst_mult_11_168 ;
wire Xd_0__inst_mult_11_169 ;
wire Xd_0__inst_mult_18_173 ;
wire Xd_0__inst_mult_18_174 ;
wire Xd_0__inst_mult_17_173 ;
wire Xd_0__inst_mult_17_174 ;
wire Xd_0__inst_mult_16_173 ;
wire Xd_0__inst_mult_16_174 ;
wire Xd_0__inst_mult_10_168 ;
wire Xd_0__inst_mult_10_169 ;
wire Xd_0__inst_mult_15_168 ;
wire Xd_0__inst_mult_15_169 ;
wire Xd_0__inst_mult_14_168 ;
wire Xd_0__inst_mult_14_169 ;
wire Xd_0__inst_mult_13_168 ;
wire Xd_0__inst_mult_13_169 ;
wire Xd_0__inst_mult_16_23_sumout ;
wire Xd_0__inst_mult_16_24 ;
wire Xd_0__inst_mult_12_168 ;
wire Xd_0__inst_mult_12_169 ;
wire Xd_0__inst_mult_15_173 ;
wire Xd_0__inst_mult_15_174 ;
wire Xd_0__inst_mult_23_28_sumout ;
wire Xd_0__inst_mult_23_29 ;
wire Xd_0__inst_mult_30_159 ;
wire Xd_0__inst_mult_30_160 ;
wire Xd_0__inst_mult_22_28_sumout ;
wire Xd_0__inst_mult_22_29 ;
wire Xd_0__inst_mult_28_154 ;
wire Xd_0__inst_mult_28_155 ;
wire Xd_0__inst_mult_0_23_sumout ;
wire Xd_0__inst_mult_0_24 ;
wire Xd_0__inst_mult_0_154 ;
wire Xd_0__inst_mult_0_155 ;
wire Xd_0__inst_mult_26_159 ;
wire Xd_0__inst_mult_26_160 ;
wire Xd_0__inst_mult_5_28_sumout ;
wire Xd_0__inst_mult_5_29 ;
wire Xd_0__inst_mult_3_154 ;
wire Xd_0__inst_mult_3_155 ;
wire Xd_0__inst_mult_16_28_sumout ;
wire Xd_0__inst_mult_16_29 ;
wire Xd_0__inst_mult_1_154 ;
wire Xd_0__inst_mult_1_155 ;
wire Xd_0__inst_mult_31_154 ;
wire Xd_0__inst_mult_31_155 ;
wire Xd_0__inst_mult_31_159 ;
wire Xd_0__inst_mult_31_160 ;
wire Xd_0__inst_mult_23_164 ;
wire Xd_0__inst_mult_23_165 ;
wire Xd_0__inst_mult_30_164 ;
wire Xd_0__inst_mult_30_165 ;
wire Xd_0__inst_mult_30_169 ;
wire Xd_0__inst_mult_30_170 ;
wire Xd_0__inst_mult_22_164 ;
wire Xd_0__inst_mult_22_165 ;
wire Xd_0__inst_mult_29_154 ;
wire Xd_0__inst_mult_29_155 ;
wire Xd_0__inst_mult_29_159 ;
wire Xd_0__inst_mult_29_160 ;
wire Xd_0__inst_mult_21_164 ;
wire Xd_0__inst_mult_21_165 ;
wire Xd_0__inst_mult_28_159 ;
wire Xd_0__inst_mult_28_160 ;
wire Xd_0__inst_mult_28_164 ;
wire Xd_0__inst_mult_28_165 ;
wire Xd_0__inst_mult_20_178 ;
wire Xd_0__inst_mult_20_179 ;
wire Xd_0__inst_mult_27_154 ;
wire Xd_0__inst_mult_27_155 ;
wire Xd_0__inst_mult_27_159 ;
wire Xd_0__inst_mult_27_160 ;
wire Xd_0__inst_mult_25_159 ;
wire Xd_0__inst_mult_25_160 ;
wire Xd_0__inst_mult_26_164 ;
wire Xd_0__inst_mult_26_165 ;
wire Xd_0__inst_mult_26_169 ;
wire Xd_0__inst_mult_26_170 ;
wire Xd_0__inst_mult_19_178 ;
wire Xd_0__inst_mult_19_179 ;
wire Xd_0__inst_mult_25_164 ;
wire Xd_0__inst_mult_25_165 ;
wire Xd_0__inst_mult_25_169 ;
wire Xd_0__inst_mult_25_170 ;
wire Xd_0__inst_mult_18_178 ;
wire Xd_0__inst_mult_18_179 ;
wire Xd_0__inst_mult_24_159 ;
wire Xd_0__inst_mult_24_160 ;
wire Xd_0__inst_mult_24_164 ;
wire Xd_0__inst_mult_24_165 ;
wire Xd_0__inst_mult_17_178 ;
wire Xd_0__inst_mult_17_179 ;
wire Xd_0__inst_mult_23_169 ;
wire Xd_0__inst_mult_23_170 ;
wire Xd_0__inst_mult_23_174 ;
wire Xd_0__inst_mult_23_175 ;
wire Xd_0__inst_mult_24_169 ;
wire Xd_0__inst_mult_24_170 ;
wire Xd_0__inst_mult_22_169 ;
wire Xd_0__inst_mult_22_170 ;
wire Xd_0__inst_mult_22_174 ;
wire Xd_0__inst_mult_22_175 ;
wire Xd_0__inst_mult_4_159 ;
wire Xd_0__inst_mult_4_160 ;
wire Xd_0__inst_mult_21_169 ;
wire Xd_0__inst_mult_21_170 ;
wire Xd_0__inst_mult_21_174 ;
wire Xd_0__inst_mult_21_175 ;
wire Xd_0__inst_mult_26_174 ;
wire Xd_0__inst_mult_26_175 ;
wire Xd_0__inst_mult_20_183 ;
wire Xd_0__inst_mult_20_184 ;
wire Xd_0__inst_mult_20_188 ;
wire Xd_0__inst_mult_20_189 ;
wire Xd_0__inst_mult_16_178 ;
wire Xd_0__inst_mult_16_179 ;
wire Xd_0__inst_mult_19_183 ;
wire Xd_0__inst_mult_19_184 ;
wire Xd_0__inst_mult_19_188 ;
wire Xd_0__inst_mult_19_189 ;
wire Xd_0__inst_mult_12_173 ;
wire Xd_0__inst_mult_12_174 ;
wire Xd_0__inst_mult_18_183 ;
wire Xd_0__inst_mult_18_184 ;
wire Xd_0__inst_mult_18_188 ;
wire Xd_0__inst_mult_18_189 ;
wire Xd_0__inst_mult_23_179 ;
wire Xd_0__inst_mult_23_180 ;
wire Xd_0__inst_mult_17_183 ;
wire Xd_0__inst_mult_17_184 ;
wire Xd_0__inst_mult_17_188 ;
wire Xd_0__inst_mult_17_189 ;
wire Xd_0__inst_mult_5_173 ;
wire Xd_0__inst_mult_5_174 ;
wire Xd_0__inst_mult_16_183 ;
wire Xd_0__inst_mult_16_184 ;
wire Xd_0__inst_mult_16_188 ;
wire Xd_0__inst_mult_16_189 ;
wire Xd_0__inst_mult_6_173 ;
wire Xd_0__inst_mult_6_174 ;
wire Xd_0__inst_mult_15_178 ;
wire Xd_0__inst_mult_15_179 ;
wire Xd_0__inst_mult_15_183 ;
wire Xd_0__inst_mult_15_184 ;
wire Xd_0__inst_mult_7_173 ;
wire Xd_0__inst_mult_7_174 ;
wire Xd_0__inst_mult_14_173 ;
wire Xd_0__inst_mult_14_174 ;
wire Xd_0__inst_mult_14_178 ;
wire Xd_0__inst_mult_14_179 ;
wire Xd_0__inst_mult_8_173 ;
wire Xd_0__inst_mult_8_174 ;
wire Xd_0__inst_mult_13_173 ;
wire Xd_0__inst_mult_13_174 ;
wire Xd_0__inst_mult_13_178 ;
wire Xd_0__inst_mult_13_179 ;
wire Xd_0__inst_mult_9_173 ;
wire Xd_0__inst_mult_9_174 ;
wire Xd_0__inst_mult_12_178 ;
wire Xd_0__inst_mult_12_179 ;
wire Xd_0__inst_mult_12_183 ;
wire Xd_0__inst_mult_12_184 ;
wire Xd_0__inst_mult_19_193 ;
wire Xd_0__inst_mult_19_194 ;
wire Xd_0__inst_mult_11_173 ;
wire Xd_0__inst_mult_11_174 ;
wire Xd_0__inst_mult_11_178 ;
wire Xd_0__inst_mult_11_179 ;
wire Xd_0__inst_mult_10_173 ;
wire Xd_0__inst_mult_10_174 ;
wire Xd_0__inst_mult_10_178 ;
wire Xd_0__inst_mult_10_179 ;
wire Xd_0__inst_mult_10_183 ;
wire Xd_0__inst_mult_10_184 ;
wire Xd_0__inst_mult_11_183 ;
wire Xd_0__inst_mult_11_184 ;
wire Xd_0__inst_mult_9_178 ;
wire Xd_0__inst_mult_9_179 ;
wire Xd_0__inst_mult_9_183 ;
wire Xd_0__inst_mult_9_184 ;
wire Xd_0__inst_mult_13_183 ;
wire Xd_0__inst_mult_13_184 ;
wire Xd_0__inst_mult_8_178 ;
wire Xd_0__inst_mult_8_179 ;
wire Xd_0__inst_mult_8_183 ;
wire Xd_0__inst_mult_8_184 ;
wire Xd_0__inst_mult_14_183 ;
wire Xd_0__inst_mult_14_184 ;
wire Xd_0__inst_mult_7_178 ;
wire Xd_0__inst_mult_7_179 ;
wire Xd_0__inst_mult_7_183 ;
wire Xd_0__inst_mult_7_184 ;
wire Xd_0__inst_mult_15_188 ;
wire Xd_0__inst_mult_15_189 ;
wire Xd_0__inst_mult_6_178 ;
wire Xd_0__inst_mult_6_179 ;
wire Xd_0__inst_mult_6_183 ;
wire Xd_0__inst_mult_6_184 ;
wire Xd_0__inst_mult_16_193 ;
wire Xd_0__inst_mult_16_194 ;
wire Xd_0__inst_mult_5_178 ;
wire Xd_0__inst_mult_5_179 ;
wire Xd_0__inst_mult_5_183 ;
wire Xd_0__inst_mult_5_184 ;
wire Xd_0__inst_mult_17_193 ;
wire Xd_0__inst_mult_17_194 ;
wire Xd_0__inst_mult_4_164 ;
wire Xd_0__inst_mult_4_165 ;
wire Xd_0__inst_mult_4_169 ;
wire Xd_0__inst_mult_4_170 ;
wire Xd_0__inst_mult_18_193 ;
wire Xd_0__inst_mult_18_194 ;
wire Xd_0__inst_mult_3_159 ;
wire Xd_0__inst_mult_3_160 ;
wire Xd_0__inst_mult_3_164 ;
wire Xd_0__inst_mult_3_165 ;
wire Xd_0__inst_mult_30_174 ;
wire Xd_0__inst_mult_30_175 ;
wire Xd_0__inst_mult_2_154 ;
wire Xd_0__inst_mult_2_155 ;
wire Xd_0__inst_mult_2_159 ;
wire Xd_0__inst_mult_2_160 ;
wire Xd_0__inst_mult_20_193 ;
wire Xd_0__inst_mult_20_194 ;
wire Xd_0__inst_mult_1_159 ;
wire Xd_0__inst_mult_1_160 ;
wire Xd_0__inst_mult_1_164 ;
wire Xd_0__inst_mult_1_165 ;
wire Xd_0__inst_mult_21_179 ;
wire Xd_0__inst_mult_21_180 ;
wire Xd_0__inst_mult_0_159 ;
wire Xd_0__inst_mult_0_160 ;
wire Xd_0__inst_mult_0_164 ;
wire Xd_0__inst_mult_0_165 ;
wire Xd_0__inst_mult_22_179 ;
wire Xd_0__inst_mult_22_180 ;
wire Xd_0__inst_mult_31_164 ;
wire Xd_0__inst_mult_31_165 ;
wire Xd_0__inst_mult_31_169 ;
wire Xd_0__inst_mult_31_170 ;
wire Xd_0__inst_mult_30_179 ;
wire Xd_0__inst_mult_30_180 ;
wire Xd_0__inst_mult_30_184 ;
wire Xd_0__inst_mult_30_185 ;
wire Xd_0__inst_mult_29_164 ;
wire Xd_0__inst_mult_29_165 ;
wire Xd_0__inst_mult_29_169 ;
wire Xd_0__inst_mult_29_170 ;
wire Xd_0__inst_mult_28_169 ;
wire Xd_0__inst_mult_28_170 ;
wire Xd_0__inst_mult_28_174 ;
wire Xd_0__inst_mult_28_175 ;
wire Xd_0__inst_mult_27_164 ;
wire Xd_0__inst_mult_27_165 ;
wire Xd_0__inst_mult_27_169 ;
wire Xd_0__inst_mult_27_170 ;
wire Xd_0__inst_mult_26_179 ;
wire Xd_0__inst_mult_26_180 ;
wire Xd_0__inst_mult_26_184 ;
wire Xd_0__inst_mult_26_185 ;
wire Xd_0__inst_mult_25_174 ;
wire Xd_0__inst_mult_25_175 ;
wire Xd_0__inst_mult_25_179 ;
wire Xd_0__inst_mult_25_180 ;
wire Xd_0__inst_mult_24_174 ;
wire Xd_0__inst_mult_24_175 ;
wire Xd_0__inst_mult_24_179 ;
wire Xd_0__inst_mult_24_180 ;
wire Xd_0__inst_mult_23_184 ;
wire Xd_0__inst_mult_23_185 ;
wire Xd_0__inst_mult_23_189 ;
wire Xd_0__inst_mult_23_190 ;
wire Xd_0__inst_mult_22_184 ;
wire Xd_0__inst_mult_22_185 ;
wire Xd_0__inst_mult_22_189 ;
wire Xd_0__inst_mult_22_190 ;
wire Xd_0__inst_mult_21_184 ;
wire Xd_0__inst_mult_21_185 ;
wire Xd_0__inst_mult_21_189 ;
wire Xd_0__inst_mult_21_190 ;
wire Xd_0__inst_mult_20_198 ;
wire Xd_0__inst_mult_20_199 ;
wire Xd_0__inst_mult_20_203 ;
wire Xd_0__inst_mult_20_204 ;
wire Xd_0__inst_mult_19_198 ;
wire Xd_0__inst_mult_19_199 ;
wire Xd_0__inst_mult_19_203 ;
wire Xd_0__inst_mult_19_204 ;
wire Xd_0__inst_mult_18_198 ;
wire Xd_0__inst_mult_18_199 ;
wire Xd_0__inst_mult_18_203 ;
wire Xd_0__inst_mult_18_204 ;
wire Xd_0__inst_mult_17_198 ;
wire Xd_0__inst_mult_17_199 ;
wire Xd_0__inst_mult_17_203 ;
wire Xd_0__inst_mult_17_204 ;
wire Xd_0__inst_mult_16_198 ;
wire Xd_0__inst_mult_16_199 ;
wire Xd_0__inst_mult_16_203 ;
wire Xd_0__inst_mult_16_204 ;
wire Xd_0__inst_mult_15_193 ;
wire Xd_0__inst_mult_15_194 ;
wire Xd_0__inst_mult_15_198 ;
wire Xd_0__inst_mult_15_199 ;
wire Xd_0__inst_mult_14_188 ;
wire Xd_0__inst_mult_14_189 ;
wire Xd_0__inst_mult_14_193 ;
wire Xd_0__inst_mult_14_194 ;
wire Xd_0__inst_mult_13_188 ;
wire Xd_0__inst_mult_13_189 ;
wire Xd_0__inst_mult_13_193 ;
wire Xd_0__inst_mult_13_194 ;
wire Xd_0__inst_mult_12_188 ;
wire Xd_0__inst_mult_12_189 ;
wire Xd_0__inst_mult_12_193 ;
wire Xd_0__inst_mult_12_194 ;
wire Xd_0__inst_mult_11_188 ;
wire Xd_0__inst_mult_11_189 ;
wire Xd_0__inst_mult_11_193 ;
wire Xd_0__inst_mult_11_194 ;
wire Xd_0__inst_mult_10_188 ;
wire Xd_0__inst_mult_10_189 ;
wire Xd_0__inst_mult_10_193 ;
wire Xd_0__inst_mult_10_194 ;
wire Xd_0__inst_mult_9_188 ;
wire Xd_0__inst_mult_9_189 ;
wire Xd_0__inst_mult_9_193 ;
wire Xd_0__inst_mult_9_194 ;
wire Xd_0__inst_mult_8_188 ;
wire Xd_0__inst_mult_8_189 ;
wire Xd_0__inst_mult_8_193 ;
wire Xd_0__inst_mult_8_194 ;
wire Xd_0__inst_mult_7_188 ;
wire Xd_0__inst_mult_7_189 ;
wire Xd_0__inst_mult_7_193 ;
wire Xd_0__inst_mult_7_194 ;
wire Xd_0__inst_mult_6_188 ;
wire Xd_0__inst_mult_6_189 ;
wire Xd_0__inst_mult_6_193 ;
wire Xd_0__inst_mult_6_194 ;
wire Xd_0__inst_mult_5_188 ;
wire Xd_0__inst_mult_5_189 ;
wire Xd_0__inst_mult_5_193 ;
wire Xd_0__inst_mult_5_194 ;
wire Xd_0__inst_mult_4_174 ;
wire Xd_0__inst_mult_4_175 ;
wire Xd_0__inst_mult_4_179 ;
wire Xd_0__inst_mult_4_180 ;
wire Xd_0__inst_mult_3_169 ;
wire Xd_0__inst_mult_3_170 ;
wire Xd_0__inst_mult_3_174 ;
wire Xd_0__inst_mult_3_175 ;
wire Xd_0__inst_mult_2_164 ;
wire Xd_0__inst_mult_2_165 ;
wire Xd_0__inst_mult_2_169 ;
wire Xd_0__inst_mult_2_170 ;
wire Xd_0__inst_mult_1_169 ;
wire Xd_0__inst_mult_1_170 ;
wire Xd_0__inst_mult_1_174 ;
wire Xd_0__inst_mult_1_175 ;
wire Xd_0__inst_mult_0_169 ;
wire Xd_0__inst_mult_0_170 ;
wire Xd_0__inst_mult_0_174 ;
wire Xd_0__inst_mult_0_175 ;
wire Xd_0__inst_mult_31_174 ;
wire Xd_0__inst_mult_31_175 ;
wire Xd_0__inst_mult_31_179 ;
wire Xd_0__inst_mult_31_180 ;
wire Xd_0__inst_mult_30_189 ;
wire Xd_0__inst_mult_30_190 ;
wire Xd_0__inst_mult_30_194 ;
wire Xd_0__inst_mult_30_195 ;
wire Xd_0__inst_mult_29_174 ;
wire Xd_0__inst_mult_29_175 ;
wire Xd_0__inst_mult_29_179 ;
wire Xd_0__inst_mult_29_180 ;
wire Xd_0__inst_mult_28_179 ;
wire Xd_0__inst_mult_28_180 ;
wire Xd_0__inst_mult_28_184 ;
wire Xd_0__inst_mult_28_185 ;
wire Xd_0__inst_mult_27_174 ;
wire Xd_0__inst_mult_27_175 ;
wire Xd_0__inst_mult_27_179 ;
wire Xd_0__inst_mult_27_180 ;
wire Xd_0__inst_mult_26_189 ;
wire Xd_0__inst_mult_26_190 ;
wire Xd_0__inst_mult_26_194 ;
wire Xd_0__inst_mult_26_195 ;
wire Xd_0__inst_mult_25_184 ;
wire Xd_0__inst_mult_25_185 ;
wire Xd_0__inst_mult_25_189 ;
wire Xd_0__inst_mult_25_190 ;
wire Xd_0__inst_mult_24_184 ;
wire Xd_0__inst_mult_24_185 ;
wire Xd_0__inst_mult_24_189 ;
wire Xd_0__inst_mult_24_190 ;
wire Xd_0__inst_mult_23_194 ;
wire Xd_0__inst_mult_23_195 ;
wire Xd_0__inst_mult_23_199 ;
wire Xd_0__inst_mult_23_200 ;
wire Xd_0__inst_mult_22_194 ;
wire Xd_0__inst_mult_22_195 ;
wire Xd_0__inst_mult_22_199 ;
wire Xd_0__inst_mult_22_200 ;
wire Xd_0__inst_mult_21_194 ;
wire Xd_0__inst_mult_21_195 ;
wire Xd_0__inst_mult_21_199 ;
wire Xd_0__inst_mult_21_200 ;
wire Xd_0__inst_mult_20_208 ;
wire Xd_0__inst_mult_20_209 ;
wire Xd_0__inst_mult_20_213 ;
wire Xd_0__inst_mult_20_214 ;
wire Xd_0__inst_mult_19_208 ;
wire Xd_0__inst_mult_19_209 ;
wire Xd_0__inst_mult_19_213 ;
wire Xd_0__inst_mult_19_214 ;
wire Xd_0__inst_mult_18_208 ;
wire Xd_0__inst_mult_18_209 ;
wire Xd_0__inst_mult_18_213 ;
wire Xd_0__inst_mult_18_214 ;
wire Xd_0__inst_mult_17_208 ;
wire Xd_0__inst_mult_17_209 ;
wire Xd_0__inst_mult_17_213 ;
wire Xd_0__inst_mult_17_214 ;
wire Xd_0__inst_mult_16_208 ;
wire Xd_0__inst_mult_16_209 ;
wire Xd_0__inst_mult_16_213 ;
wire Xd_0__inst_mult_16_214 ;
wire Xd_0__inst_mult_15_203 ;
wire Xd_0__inst_mult_15_204 ;
wire Xd_0__inst_mult_15_208 ;
wire Xd_0__inst_mult_15_209 ;
wire Xd_0__inst_mult_14_198 ;
wire Xd_0__inst_mult_14_199 ;
wire Xd_0__inst_mult_14_203 ;
wire Xd_0__inst_mult_14_204 ;
wire Xd_0__inst_mult_13_198 ;
wire Xd_0__inst_mult_13_199 ;
wire Xd_0__inst_mult_13_203 ;
wire Xd_0__inst_mult_13_204 ;
wire Xd_0__inst_mult_12_198 ;
wire Xd_0__inst_mult_12_199 ;
wire Xd_0__inst_mult_12_203 ;
wire Xd_0__inst_mult_12_204 ;
wire Xd_0__inst_mult_11_198 ;
wire Xd_0__inst_mult_11_199 ;
wire Xd_0__inst_mult_11_203 ;
wire Xd_0__inst_mult_11_204 ;
wire Xd_0__inst_mult_10_198 ;
wire Xd_0__inst_mult_10_199 ;
wire Xd_0__inst_mult_10_203 ;
wire Xd_0__inst_mult_10_204 ;
wire Xd_0__inst_mult_9_198 ;
wire Xd_0__inst_mult_9_199 ;
wire Xd_0__inst_mult_9_203 ;
wire Xd_0__inst_mult_9_204 ;
wire Xd_0__inst_mult_8_198 ;
wire Xd_0__inst_mult_8_199 ;
wire Xd_0__inst_mult_8_203 ;
wire Xd_0__inst_mult_8_204 ;
wire Xd_0__inst_mult_7_198 ;
wire Xd_0__inst_mult_7_199 ;
wire Xd_0__inst_mult_7_203 ;
wire Xd_0__inst_mult_7_204 ;
wire Xd_0__inst_mult_6_198 ;
wire Xd_0__inst_mult_6_199 ;
wire Xd_0__inst_mult_6_203 ;
wire Xd_0__inst_mult_6_204 ;
wire Xd_0__inst_mult_5_198 ;
wire Xd_0__inst_mult_5_199 ;
wire Xd_0__inst_mult_5_203 ;
wire Xd_0__inst_mult_5_204 ;
wire Xd_0__inst_mult_4_184 ;
wire Xd_0__inst_mult_4_185 ;
wire Xd_0__inst_mult_4_189 ;
wire Xd_0__inst_mult_4_190 ;
wire Xd_0__inst_mult_3_179 ;
wire Xd_0__inst_mult_3_180 ;
wire Xd_0__inst_mult_3_184 ;
wire Xd_0__inst_mult_3_185 ;
wire Xd_0__inst_mult_2_174 ;
wire Xd_0__inst_mult_2_175 ;
wire Xd_0__inst_mult_2_179 ;
wire Xd_0__inst_mult_2_180 ;
wire Xd_0__inst_mult_1_179 ;
wire Xd_0__inst_mult_1_180 ;
wire Xd_0__inst_mult_1_184 ;
wire Xd_0__inst_mult_1_185 ;
wire Xd_0__inst_mult_0_179 ;
wire Xd_0__inst_mult_0_180 ;
wire Xd_0__inst_mult_0_184 ;
wire Xd_0__inst_mult_0_185 ;
wire Xd_0__inst_mult_31_184 ;
wire Xd_0__inst_mult_31_185 ;
wire Xd_0__inst_mult_31_189 ;
wire Xd_0__inst_mult_31_190 ;
wire Xd_0__inst_mult_30_199 ;
wire Xd_0__inst_mult_30_200 ;
wire Xd_0__inst_mult_30_204 ;
wire Xd_0__inst_mult_30_205 ;
wire Xd_0__inst_mult_29_184 ;
wire Xd_0__inst_mult_29_185 ;
wire Xd_0__inst_mult_29_189 ;
wire Xd_0__inst_mult_29_190 ;
wire Xd_0__inst_mult_28_189 ;
wire Xd_0__inst_mult_28_190 ;
wire Xd_0__inst_mult_28_194 ;
wire Xd_0__inst_mult_28_195 ;
wire Xd_0__inst_mult_27_184 ;
wire Xd_0__inst_mult_27_185 ;
wire Xd_0__inst_mult_27_189 ;
wire Xd_0__inst_mult_27_190 ;
wire Xd_0__inst_mult_26_199 ;
wire Xd_0__inst_mult_26_200 ;
wire Xd_0__inst_mult_26_204 ;
wire Xd_0__inst_mult_26_205 ;
wire Xd_0__inst_mult_25_194 ;
wire Xd_0__inst_mult_25_195 ;
wire Xd_0__inst_mult_25_199 ;
wire Xd_0__inst_mult_25_200 ;
wire Xd_0__inst_mult_24_194 ;
wire Xd_0__inst_mult_24_195 ;
wire Xd_0__inst_mult_24_199 ;
wire Xd_0__inst_mult_24_200 ;
wire Xd_0__inst_mult_23_204 ;
wire Xd_0__inst_mult_23_205 ;
wire Xd_0__inst_mult_23_209 ;
wire Xd_0__inst_mult_23_210 ;
wire Xd_0__inst_mult_22_204 ;
wire Xd_0__inst_mult_22_205 ;
wire Xd_0__inst_mult_22_209 ;
wire Xd_0__inst_mult_22_210 ;
wire Xd_0__inst_mult_21_204 ;
wire Xd_0__inst_mult_21_205 ;
wire Xd_0__inst_mult_21_209 ;
wire Xd_0__inst_mult_21_210 ;
wire Xd_0__inst_mult_20_218 ;
wire Xd_0__inst_mult_20_219 ;
wire Xd_0__inst_mult_20_223 ;
wire Xd_0__inst_mult_20_224 ;
wire Xd_0__inst_mult_19_218 ;
wire Xd_0__inst_mult_19_219 ;
wire Xd_0__inst_mult_19_223 ;
wire Xd_0__inst_mult_19_224 ;
wire Xd_0__inst_mult_18_218 ;
wire Xd_0__inst_mult_18_219 ;
wire Xd_0__inst_mult_18_223 ;
wire Xd_0__inst_mult_18_224 ;
wire Xd_0__inst_mult_17_218 ;
wire Xd_0__inst_mult_17_219 ;
wire Xd_0__inst_mult_17_223 ;
wire Xd_0__inst_mult_17_224 ;
wire Xd_0__inst_mult_16_218 ;
wire Xd_0__inst_mult_16_219 ;
wire Xd_0__inst_mult_16_223 ;
wire Xd_0__inst_mult_16_224 ;
wire Xd_0__inst_mult_15_213 ;
wire Xd_0__inst_mult_15_214 ;
wire Xd_0__inst_mult_15_218 ;
wire Xd_0__inst_mult_15_219 ;
wire Xd_0__inst_mult_14_208 ;
wire Xd_0__inst_mult_14_209 ;
wire Xd_0__inst_mult_14_213 ;
wire Xd_0__inst_mult_14_214 ;
wire Xd_0__inst_mult_13_208 ;
wire Xd_0__inst_mult_13_209 ;
wire Xd_0__inst_mult_13_213 ;
wire Xd_0__inst_mult_13_214 ;
wire Xd_0__inst_mult_12_208 ;
wire Xd_0__inst_mult_12_209 ;
wire Xd_0__inst_mult_12_213 ;
wire Xd_0__inst_mult_12_214 ;
wire Xd_0__inst_mult_11_208 ;
wire Xd_0__inst_mult_11_209 ;
wire Xd_0__inst_mult_11_213 ;
wire Xd_0__inst_mult_11_214 ;
wire Xd_0__inst_mult_10_208 ;
wire Xd_0__inst_mult_10_209 ;
wire Xd_0__inst_mult_10_213 ;
wire Xd_0__inst_mult_10_214 ;
wire Xd_0__inst_mult_9_208 ;
wire Xd_0__inst_mult_9_209 ;
wire Xd_0__inst_mult_9_213 ;
wire Xd_0__inst_mult_9_214 ;
wire Xd_0__inst_mult_8_208 ;
wire Xd_0__inst_mult_8_209 ;
wire Xd_0__inst_mult_8_213 ;
wire Xd_0__inst_mult_8_214 ;
wire Xd_0__inst_mult_7_208 ;
wire Xd_0__inst_mult_7_209 ;
wire Xd_0__inst_mult_7_213 ;
wire Xd_0__inst_mult_7_214 ;
wire Xd_0__inst_mult_6_208 ;
wire Xd_0__inst_mult_6_209 ;
wire Xd_0__inst_mult_6_213 ;
wire Xd_0__inst_mult_6_214 ;
wire Xd_0__inst_mult_5_208 ;
wire Xd_0__inst_mult_5_209 ;
wire Xd_0__inst_mult_5_213 ;
wire Xd_0__inst_mult_5_214 ;
wire Xd_0__inst_mult_4_194 ;
wire Xd_0__inst_mult_4_195 ;
wire Xd_0__inst_mult_4_199 ;
wire Xd_0__inst_mult_4_200 ;
wire Xd_0__inst_mult_3_189 ;
wire Xd_0__inst_mult_3_190 ;
wire Xd_0__inst_mult_3_194 ;
wire Xd_0__inst_mult_3_195 ;
wire Xd_0__inst_mult_2_184 ;
wire Xd_0__inst_mult_2_185 ;
wire Xd_0__inst_mult_2_189 ;
wire Xd_0__inst_mult_2_190 ;
wire Xd_0__inst_mult_1_189 ;
wire Xd_0__inst_mult_1_190 ;
wire Xd_0__inst_mult_1_194 ;
wire Xd_0__inst_mult_1_195 ;
wire Xd_0__inst_mult_0_189 ;
wire Xd_0__inst_mult_0_190 ;
wire Xd_0__inst_mult_0_194 ;
wire Xd_0__inst_mult_0_195 ;
wire Xd_0__inst_mult_31_194 ;
wire Xd_0__inst_mult_31_195 ;
wire Xd_0__inst_mult_31_199 ;
wire Xd_0__inst_mult_31_200 ;
wire Xd_0__inst_mult_30_209 ;
wire Xd_0__inst_mult_30_210 ;
wire Xd_0__inst_mult_30_214 ;
wire Xd_0__inst_mult_30_215 ;
wire Xd_0__inst_mult_29_194 ;
wire Xd_0__inst_mult_29_195 ;
wire Xd_0__inst_mult_29_199 ;
wire Xd_0__inst_mult_29_200 ;
wire Xd_0__inst_mult_28_199 ;
wire Xd_0__inst_mult_28_200 ;
wire Xd_0__inst_mult_28_204 ;
wire Xd_0__inst_mult_28_205 ;
wire Xd_0__inst_mult_27_194 ;
wire Xd_0__inst_mult_27_195 ;
wire Xd_0__inst_mult_27_199 ;
wire Xd_0__inst_mult_27_200 ;
wire Xd_0__inst_mult_26_209 ;
wire Xd_0__inst_mult_26_210 ;
wire Xd_0__inst_mult_26_214 ;
wire Xd_0__inst_mult_26_215 ;
wire Xd_0__inst_mult_25_204 ;
wire Xd_0__inst_mult_25_205 ;
wire Xd_0__inst_mult_25_209 ;
wire Xd_0__inst_mult_25_210 ;
wire Xd_0__inst_mult_24_204 ;
wire Xd_0__inst_mult_24_205 ;
wire Xd_0__inst_mult_24_209 ;
wire Xd_0__inst_mult_24_210 ;
wire Xd_0__inst_mult_23_214 ;
wire Xd_0__inst_mult_23_215 ;
wire Xd_0__inst_mult_23_219 ;
wire Xd_0__inst_mult_23_220 ;
wire Xd_0__inst_mult_22_214 ;
wire Xd_0__inst_mult_22_215 ;
wire Xd_0__inst_mult_22_219 ;
wire Xd_0__inst_mult_22_220 ;
wire Xd_0__inst_mult_21_214 ;
wire Xd_0__inst_mult_21_215 ;
wire Xd_0__inst_mult_21_219 ;
wire Xd_0__inst_mult_21_220 ;
wire Xd_0__inst_mult_20_228 ;
wire Xd_0__inst_mult_20_229 ;
wire Xd_0__inst_mult_20_233 ;
wire Xd_0__inst_mult_20_234 ;
wire Xd_0__inst_mult_19_228 ;
wire Xd_0__inst_mult_19_229 ;
wire Xd_0__inst_mult_19_233 ;
wire Xd_0__inst_mult_19_234 ;
wire Xd_0__inst_mult_18_228 ;
wire Xd_0__inst_mult_18_229 ;
wire Xd_0__inst_mult_18_233 ;
wire Xd_0__inst_mult_18_234 ;
wire Xd_0__inst_mult_17_228 ;
wire Xd_0__inst_mult_17_229 ;
wire Xd_0__inst_mult_17_233 ;
wire Xd_0__inst_mult_17_234 ;
wire Xd_0__inst_mult_16_228 ;
wire Xd_0__inst_mult_16_229 ;
wire Xd_0__inst_mult_16_233 ;
wire Xd_0__inst_mult_16_234 ;
wire Xd_0__inst_mult_15_223 ;
wire Xd_0__inst_mult_15_224 ;
wire Xd_0__inst_mult_15_228 ;
wire Xd_0__inst_mult_15_229 ;
wire Xd_0__inst_mult_14_218 ;
wire Xd_0__inst_mult_14_219 ;
wire Xd_0__inst_mult_14_223 ;
wire Xd_0__inst_mult_14_224 ;
wire Xd_0__inst_mult_13_218 ;
wire Xd_0__inst_mult_13_219 ;
wire Xd_0__inst_mult_13_223 ;
wire Xd_0__inst_mult_13_224 ;
wire Xd_0__inst_mult_12_218 ;
wire Xd_0__inst_mult_12_219 ;
wire Xd_0__inst_mult_12_223 ;
wire Xd_0__inst_mult_12_224 ;
wire Xd_0__inst_mult_11_218 ;
wire Xd_0__inst_mult_11_219 ;
wire Xd_0__inst_mult_11_223 ;
wire Xd_0__inst_mult_11_224 ;
wire Xd_0__inst_mult_10_218 ;
wire Xd_0__inst_mult_10_219 ;
wire Xd_0__inst_mult_10_223 ;
wire Xd_0__inst_mult_10_224 ;
wire Xd_0__inst_mult_9_218 ;
wire Xd_0__inst_mult_9_219 ;
wire Xd_0__inst_mult_9_223 ;
wire Xd_0__inst_mult_9_224 ;
wire Xd_0__inst_mult_8_218 ;
wire Xd_0__inst_mult_8_219 ;
wire Xd_0__inst_mult_8_223 ;
wire Xd_0__inst_mult_8_224 ;
wire Xd_0__inst_mult_7_218 ;
wire Xd_0__inst_mult_7_219 ;
wire Xd_0__inst_mult_7_223 ;
wire Xd_0__inst_mult_7_224 ;
wire Xd_0__inst_mult_6_218 ;
wire Xd_0__inst_mult_6_219 ;
wire Xd_0__inst_mult_6_223 ;
wire Xd_0__inst_mult_6_224 ;
wire Xd_0__inst_mult_5_218 ;
wire Xd_0__inst_mult_5_219 ;
wire Xd_0__inst_mult_5_223 ;
wire Xd_0__inst_mult_5_224 ;
wire Xd_0__inst_mult_4_204 ;
wire Xd_0__inst_mult_4_205 ;
wire Xd_0__inst_mult_4_209 ;
wire Xd_0__inst_mult_4_210 ;
wire Xd_0__inst_mult_3_199 ;
wire Xd_0__inst_mult_3_200 ;
wire Xd_0__inst_mult_3_204 ;
wire Xd_0__inst_mult_3_205 ;
wire Xd_0__inst_mult_2_194 ;
wire Xd_0__inst_mult_2_195 ;
wire Xd_0__inst_mult_2_199 ;
wire Xd_0__inst_mult_2_200 ;
wire Xd_0__inst_mult_1_199 ;
wire Xd_0__inst_mult_1_200 ;
wire Xd_0__inst_mult_1_204 ;
wire Xd_0__inst_mult_1_205 ;
wire Xd_0__inst_mult_0_199 ;
wire Xd_0__inst_mult_0_200 ;
wire Xd_0__inst_mult_0_204 ;
wire Xd_0__inst_mult_0_205 ;
wire Xd_0__inst_mult_31_204 ;
wire Xd_0__inst_mult_31_205 ;
wire Xd_0__inst_mult_31_209 ;
wire Xd_0__inst_mult_31_210 ;
wire Xd_0__inst_mult_30_219 ;
wire Xd_0__inst_mult_30_220 ;
wire Xd_0__inst_mult_30_224 ;
wire Xd_0__inst_mult_30_225 ;
wire Xd_0__inst_mult_29_204 ;
wire Xd_0__inst_mult_29_205 ;
wire Xd_0__inst_mult_29_209 ;
wire Xd_0__inst_mult_29_210 ;
wire Xd_0__inst_mult_28_209 ;
wire Xd_0__inst_mult_28_210 ;
wire Xd_0__inst_mult_28_214 ;
wire Xd_0__inst_mult_28_215 ;
wire Xd_0__inst_mult_27_204 ;
wire Xd_0__inst_mult_27_205 ;
wire Xd_0__inst_mult_27_209 ;
wire Xd_0__inst_mult_27_210 ;
wire Xd_0__inst_mult_26_219 ;
wire Xd_0__inst_mult_26_220 ;
wire Xd_0__inst_mult_26_224 ;
wire Xd_0__inst_mult_26_225 ;
wire Xd_0__inst_mult_25_214 ;
wire Xd_0__inst_mult_25_215 ;
wire Xd_0__inst_mult_25_219 ;
wire Xd_0__inst_mult_25_220 ;
wire Xd_0__inst_mult_24_214 ;
wire Xd_0__inst_mult_24_215 ;
wire Xd_0__inst_mult_24_219 ;
wire Xd_0__inst_mult_24_220 ;
wire Xd_0__inst_mult_23_224 ;
wire Xd_0__inst_mult_23_225 ;
wire Xd_0__inst_mult_23_229 ;
wire Xd_0__inst_mult_23_230 ;
wire Xd_0__inst_mult_22_224 ;
wire Xd_0__inst_mult_22_225 ;
wire Xd_0__inst_mult_22_229 ;
wire Xd_0__inst_mult_22_230 ;
wire Xd_0__inst_mult_21_224 ;
wire Xd_0__inst_mult_21_225 ;
wire Xd_0__inst_mult_21_229 ;
wire Xd_0__inst_mult_21_230 ;
wire Xd_0__inst_mult_20_238 ;
wire Xd_0__inst_mult_20_239 ;
wire Xd_0__inst_mult_20_243 ;
wire Xd_0__inst_mult_20_244 ;
wire Xd_0__inst_mult_19_238 ;
wire Xd_0__inst_mult_19_239 ;
wire Xd_0__inst_mult_19_243 ;
wire Xd_0__inst_mult_19_244 ;
wire Xd_0__inst_mult_18_238 ;
wire Xd_0__inst_mult_18_239 ;
wire Xd_0__inst_mult_18_243 ;
wire Xd_0__inst_mult_18_244 ;
wire Xd_0__inst_mult_17_238 ;
wire Xd_0__inst_mult_17_239 ;
wire Xd_0__inst_mult_17_243 ;
wire Xd_0__inst_mult_17_244 ;
wire Xd_0__inst_mult_16_238 ;
wire Xd_0__inst_mult_16_239 ;
wire Xd_0__inst_mult_16_243 ;
wire Xd_0__inst_mult_16_244 ;
wire Xd_0__inst_mult_15_233 ;
wire Xd_0__inst_mult_15_234 ;
wire Xd_0__inst_mult_15_238 ;
wire Xd_0__inst_mult_15_239 ;
wire Xd_0__inst_mult_14_228 ;
wire Xd_0__inst_mult_14_229 ;
wire Xd_0__inst_mult_14_233 ;
wire Xd_0__inst_mult_14_234 ;
wire Xd_0__inst_mult_13_228 ;
wire Xd_0__inst_mult_13_229 ;
wire Xd_0__inst_mult_13_233 ;
wire Xd_0__inst_mult_13_234 ;
wire Xd_0__inst_mult_12_228 ;
wire Xd_0__inst_mult_12_229 ;
wire Xd_0__inst_mult_12_233 ;
wire Xd_0__inst_mult_12_234 ;
wire Xd_0__inst_mult_11_228 ;
wire Xd_0__inst_mult_11_229 ;
wire Xd_0__inst_mult_11_233 ;
wire Xd_0__inst_mult_11_234 ;
wire Xd_0__inst_mult_10_228 ;
wire Xd_0__inst_mult_10_229 ;
wire Xd_0__inst_mult_10_233 ;
wire Xd_0__inst_mult_10_234 ;
wire Xd_0__inst_mult_9_228 ;
wire Xd_0__inst_mult_9_229 ;
wire Xd_0__inst_mult_9_233 ;
wire Xd_0__inst_mult_9_234 ;
wire Xd_0__inst_mult_8_228 ;
wire Xd_0__inst_mult_8_229 ;
wire Xd_0__inst_mult_8_233 ;
wire Xd_0__inst_mult_8_234 ;
wire Xd_0__inst_mult_7_228 ;
wire Xd_0__inst_mult_7_229 ;
wire Xd_0__inst_mult_7_233 ;
wire Xd_0__inst_mult_7_234 ;
wire Xd_0__inst_mult_6_228 ;
wire Xd_0__inst_mult_6_229 ;
wire Xd_0__inst_mult_6_233 ;
wire Xd_0__inst_mult_6_234 ;
wire Xd_0__inst_mult_5_228 ;
wire Xd_0__inst_mult_5_229 ;
wire Xd_0__inst_mult_5_233 ;
wire Xd_0__inst_mult_5_234 ;
wire Xd_0__inst_mult_4_214 ;
wire Xd_0__inst_mult_4_215 ;
wire Xd_0__inst_mult_4_219 ;
wire Xd_0__inst_mult_4_220 ;
wire Xd_0__inst_mult_3_209 ;
wire Xd_0__inst_mult_3_210 ;
wire Xd_0__inst_mult_3_214 ;
wire Xd_0__inst_mult_3_215 ;
wire Xd_0__inst_mult_2_204 ;
wire Xd_0__inst_mult_2_205 ;
wire Xd_0__inst_mult_2_209 ;
wire Xd_0__inst_mult_2_210 ;
wire Xd_0__inst_mult_1_209 ;
wire Xd_0__inst_mult_1_210 ;
wire Xd_0__inst_mult_1_214 ;
wire Xd_0__inst_mult_1_215 ;
wire Xd_0__inst_mult_0_209 ;
wire Xd_0__inst_mult_0_210 ;
wire Xd_0__inst_mult_0_214 ;
wire Xd_0__inst_mult_0_215 ;
wire Xd_0__inst_mult_31_214 ;
wire Xd_0__inst_mult_31_219 ;
wire Xd_0__inst_mult_31_220 ;
wire Xd_0__inst_mult_30_229 ;
wire Xd_0__inst_mult_30_230 ;
wire Xd_0__inst_mult_30_234 ;
wire Xd_0__inst_mult_30_235 ;
wire Xd_0__inst_mult_29_214 ;
wire Xd_0__inst_mult_29_219 ;
wire Xd_0__inst_mult_29_220 ;
wire Xd_0__inst_mult_28_219 ;
wire Xd_0__inst_mult_28_220 ;
wire Xd_0__inst_mult_28_224 ;
wire Xd_0__inst_mult_28_225 ;
wire Xd_0__inst_mult_27_214 ;
wire Xd_0__inst_mult_27_219 ;
wire Xd_0__inst_mult_27_220 ;
wire Xd_0__inst_mult_26_229 ;
wire Xd_0__inst_mult_26_230 ;
wire Xd_0__inst_mult_26_234 ;
wire Xd_0__inst_mult_26_235 ;
wire Xd_0__inst_mult_25_224 ;
wire Xd_0__inst_mult_25_229 ;
wire Xd_0__inst_mult_25_230 ;
wire Xd_0__inst_mult_24_224 ;
wire Xd_0__inst_mult_24_225 ;
wire Xd_0__inst_mult_24_229 ;
wire Xd_0__inst_mult_24_230 ;
wire Xd_0__inst_mult_23_234 ;
wire Xd_0__inst_mult_23_235 ;
wire Xd_0__inst_mult_23_239 ;
wire Xd_0__inst_mult_23_240 ;
wire Xd_0__inst_mult_22_234 ;
wire Xd_0__inst_mult_22_239 ;
wire Xd_0__inst_mult_22_240 ;
wire Xd_0__inst_mult_21_234 ;
wire Xd_0__inst_mult_21_235 ;
wire Xd_0__inst_mult_21_239 ;
wire Xd_0__inst_mult_21_240 ;
wire Xd_0__inst_mult_20_248 ;
wire Xd_0__inst_mult_20_253 ;
wire Xd_0__inst_mult_20_254 ;
wire Xd_0__inst_mult_19_248 ;
wire Xd_0__inst_mult_19_249 ;
wire Xd_0__inst_mult_19_253 ;
wire Xd_0__inst_mult_19_254 ;
wire Xd_0__inst_mult_18_248 ;
wire Xd_0__inst_mult_18_253 ;
wire Xd_0__inst_mult_18_254 ;
wire Xd_0__inst_mult_17_248 ;
wire Xd_0__inst_mult_17_253 ;
wire Xd_0__inst_mult_17_254 ;
wire Xd_0__inst_mult_16_248 ;
wire Xd_0__inst_mult_16_249 ;
wire Xd_0__inst_mult_16_253 ;
wire Xd_0__inst_mult_16_254 ;
wire Xd_0__inst_mult_15_243 ;
wire Xd_0__inst_mult_15_248 ;
wire Xd_0__inst_mult_15_249 ;
wire Xd_0__inst_mult_14_238 ;
wire Xd_0__inst_mult_14_239 ;
wire Xd_0__inst_mult_14_243 ;
wire Xd_0__inst_mult_14_244 ;
wire Xd_0__inst_mult_13_238 ;
wire Xd_0__inst_mult_13_243 ;
wire Xd_0__inst_mult_13_244 ;
wire Xd_0__inst_mult_12_238 ;
wire Xd_0__inst_mult_12_239 ;
wire Xd_0__inst_mult_12_243 ;
wire Xd_0__inst_mult_12_244 ;
wire Xd_0__inst_mult_11_238 ;
wire Xd_0__inst_mult_11_243 ;
wire Xd_0__inst_mult_11_244 ;
wire Xd_0__inst_mult_10_238 ;
wire Xd_0__inst_mult_10_239 ;
wire Xd_0__inst_mult_10_243 ;
wire Xd_0__inst_mult_10_244 ;
wire Xd_0__inst_mult_9_238 ;
wire Xd_0__inst_mult_9_243 ;
wire Xd_0__inst_mult_9_244 ;
wire Xd_0__inst_mult_8_238 ;
wire Xd_0__inst_mult_8_239 ;
wire Xd_0__inst_mult_8_243 ;
wire Xd_0__inst_mult_8_244 ;
wire Xd_0__inst_mult_7_238 ;
wire Xd_0__inst_mult_7_243 ;
wire Xd_0__inst_mult_7_244 ;
wire Xd_0__inst_mult_6_238 ;
wire Xd_0__inst_mult_6_239 ;
wire Xd_0__inst_mult_6_243 ;
wire Xd_0__inst_mult_6_244 ;
wire Xd_0__inst_mult_5_238 ;
wire Xd_0__inst_mult_5_243 ;
wire Xd_0__inst_mult_5_244 ;
wire Xd_0__inst_mult_4_224 ;
wire Xd_0__inst_mult_4_225 ;
wire Xd_0__inst_mult_4_229 ;
wire Xd_0__inst_mult_4_230 ;
wire Xd_0__inst_mult_3_219 ;
wire Xd_0__inst_mult_3_224 ;
wire Xd_0__inst_mult_3_225 ;
wire Xd_0__inst_mult_2_214 ;
wire Xd_0__inst_mult_2_215 ;
wire Xd_0__inst_mult_2_219 ;
wire Xd_0__inst_mult_2_220 ;
wire Xd_0__inst_mult_1_219 ;
wire Xd_0__inst_mult_1_224 ;
wire Xd_0__inst_mult_1_225 ;
wire Xd_0__inst_mult_0_219 ;
wire Xd_0__inst_mult_0_220 ;
wire Xd_0__inst_mult_0_224 ;
wire Xd_0__inst_mult_0_225 ;
wire Xd_0__inst_mult_31_224 ;
wire Xd_0__inst_mult_31_225 ;
wire Xd_0__inst_mult_31_28_sumout ;
wire Xd_0__inst_mult_31_29 ;
wire Xd_0__inst_mult_30_239 ;
wire Xd_0__inst_mult_30_240 ;
wire Xd_0__inst_mult_30_28_sumout ;
wire Xd_0__inst_mult_30_29 ;
wire Xd_0__inst_mult_29_224 ;
wire Xd_0__inst_mult_29_225 ;
wire Xd_0__inst_mult_29_28_sumout ;
wire Xd_0__inst_mult_29_29 ;
wire Xd_0__inst_mult_28_229 ;
wire Xd_0__inst_mult_28_230 ;
wire Xd_0__inst_mult_28_28_sumout ;
wire Xd_0__inst_mult_28_29 ;
wire Xd_0__inst_mult_27_224 ;
wire Xd_0__inst_mult_27_225 ;
wire Xd_0__inst_mult_27_28_sumout ;
wire Xd_0__inst_mult_27_29 ;
wire Xd_0__inst_mult_26_239 ;
wire Xd_0__inst_mult_26_240 ;
wire Xd_0__inst_mult_26_28_sumout ;
wire Xd_0__inst_mult_25_234 ;
wire Xd_0__inst_mult_25_235 ;
wire Xd_0__inst_mult_25_28_sumout ;
wire Xd_0__inst_mult_25_29 ;
wire Xd_0__inst_mult_24_234 ;
wire Xd_0__inst_mult_24_235 ;
wire Xd_0__inst_mult_24_28_sumout ;
wire Xd_0__inst_mult_24_29 ;
wire Xd_0__inst_mult_23_244 ;
wire Xd_0__inst_mult_23_245 ;
wire Xd_0__inst_mult_23_33_sumout ;
wire Xd_0__inst_mult_23_34 ;
wire Xd_0__inst_mult_22_244 ;
wire Xd_0__inst_mult_22_245 ;
wire Xd_0__inst_mult_22_33_sumout ;
wire Xd_0__inst_mult_22_34 ;
wire Xd_0__inst_mult_21_244 ;
wire Xd_0__inst_mult_21_245 ;
wire Xd_0__inst_mult_21_28_sumout ;
wire Xd_0__inst_mult_21_29 ;
wire Xd_0__inst_mult_20_258 ;
wire Xd_0__inst_mult_20_259 ;
wire Xd_0__inst_mult_20_23_sumout ;
wire Xd_0__inst_mult_20_24 ;
wire Xd_0__inst_mult_19_258 ;
wire Xd_0__inst_mult_19_259 ;
wire Xd_0__inst_mult_19_23_sumout ;
wire Xd_0__inst_mult_19_24 ;
wire Xd_0__inst_mult_18_258 ;
wire Xd_0__inst_mult_18_259 ;
wire Xd_0__inst_mult_18_23_sumout ;
wire Xd_0__inst_mult_18_24 ;
wire Xd_0__inst_mult_17_258 ;
wire Xd_0__inst_mult_17_259 ;
wire Xd_0__inst_mult_17_23_sumout ;
wire Xd_0__inst_mult_17_24 ;
wire Xd_0__inst_mult_16_258 ;
wire Xd_0__inst_mult_16_259 ;
wire Xd_0__inst_mult_15_253 ;
wire Xd_0__inst_mult_15_254 ;
wire Xd_0__inst_mult_15_23_sumout ;
wire Xd_0__inst_mult_15_24 ;
wire Xd_0__inst_mult_14_248 ;
wire Xd_0__inst_mult_14_249 ;
wire Xd_0__inst_mult_14_28_sumout ;
wire Xd_0__inst_mult_14_29 ;
wire Xd_0__inst_mult_13_248 ;
wire Xd_0__inst_mult_13_249 ;
wire Xd_0__inst_mult_13_28_sumout ;
wire Xd_0__inst_mult_13_29 ;
wire Xd_0__inst_mult_12_248 ;
wire Xd_0__inst_mult_12_249 ;
wire Xd_0__inst_mult_12_28_sumout ;
wire Xd_0__inst_mult_12_29 ;
wire Xd_0__inst_mult_11_248 ;
wire Xd_0__inst_mult_11_249 ;
wire Xd_0__inst_mult_11_28_sumout ;
wire Xd_0__inst_mult_11_29 ;
wire Xd_0__inst_mult_10_248 ;
wire Xd_0__inst_mult_10_249 ;
wire Xd_0__inst_mult_10_33_sumout ;
wire Xd_0__inst_mult_10_34 ;
wire Xd_0__inst_mult_9_248 ;
wire Xd_0__inst_mult_9_249 ;
wire Xd_0__inst_mult_9_28_sumout ;
wire Xd_0__inst_mult_9_29 ;
wire Xd_0__inst_mult_8_248 ;
wire Xd_0__inst_mult_8_249 ;
wire Xd_0__inst_mult_8_28_sumout ;
wire Xd_0__inst_mult_8_29 ;
wire Xd_0__inst_mult_7_248 ;
wire Xd_0__inst_mult_7_249 ;
wire Xd_0__inst_mult_7_28_sumout ;
wire Xd_0__inst_mult_7_29 ;
wire Xd_0__inst_mult_6_248 ;
wire Xd_0__inst_mult_6_249 ;
wire Xd_0__inst_mult_6_28_sumout ;
wire Xd_0__inst_mult_6_29 ;
wire Xd_0__inst_mult_5_248 ;
wire Xd_0__inst_mult_5_249 ;
wire Xd_0__inst_mult_5_33_sumout ;
wire Xd_0__inst_mult_5_34 ;
wire Xd_0__inst_mult_4_234 ;
wire Xd_0__inst_mult_4_235 ;
wire Xd_0__inst_mult_4_28_sumout ;
wire Xd_0__inst_mult_4_29 ;
wire Xd_0__inst_mult_3_229 ;
wire Xd_0__inst_mult_3_230 ;
wire Xd_0__inst_mult_3_28_sumout ;
wire Xd_0__inst_mult_3_29 ;
wire Xd_0__inst_mult_2_224 ;
wire Xd_0__inst_mult_2_225 ;
wire Xd_0__inst_mult_2_28_sumout ;
wire Xd_0__inst_mult_2_29 ;
wire Xd_0__inst_mult_1_229 ;
wire Xd_0__inst_mult_1_230 ;
wire Xd_0__inst_mult_1_28_sumout ;
wire Xd_0__inst_mult_1_29 ;
wire Xd_0__inst_mult_0_229 ;
wire Xd_0__inst_mult_0_230 ;
wire Xd_0__inst_mult_0_28_sumout ;
wire Xd_0__inst_mult_0_29 ;
wire Xd_0__inst_mult_31_229 ;
wire Xd_0__inst_mult_31_230 ;
wire Xd_0__inst_mult_30_244 ;
wire Xd_0__inst_mult_30_245 ;
wire Xd_0__inst_mult_29_229 ;
wire Xd_0__inst_mult_29_230 ;
wire Xd_0__inst_mult_28_234 ;
wire Xd_0__inst_mult_28_235 ;
wire Xd_0__inst_mult_27_229 ;
wire Xd_0__inst_mult_27_230 ;
wire Xd_0__inst_mult_26_244 ;
wire Xd_0__inst_mult_26_245 ;
wire Xd_0__inst_mult_25_239 ;
wire Xd_0__inst_mult_25_240 ;
wire Xd_0__inst_mult_24_239 ;
wire Xd_0__inst_mult_24_240 ;
wire Xd_0__inst_mult_23_249 ;
wire Xd_0__inst_mult_23_250 ;
wire Xd_0__inst_mult_22_249 ;
wire Xd_0__inst_mult_22_250 ;
wire Xd_0__inst_mult_21_249 ;
wire Xd_0__inst_mult_21_250 ;
wire Xd_0__inst_mult_20_263 ;
wire Xd_0__inst_mult_20_264 ;
wire Xd_0__inst_mult_20_28_sumout ;
wire Xd_0__inst_mult_20_29 ;
wire Xd_0__inst_mult_19_263 ;
wire Xd_0__inst_mult_19_264 ;
wire Xd_0__inst_mult_19_28_sumout ;
wire Xd_0__inst_mult_19_29 ;
wire Xd_0__inst_mult_18_263 ;
wire Xd_0__inst_mult_18_264 ;
wire Xd_0__inst_mult_18_28_sumout ;
wire Xd_0__inst_mult_18_29 ;
wire Xd_0__inst_mult_17_263 ;
wire Xd_0__inst_mult_17_264 ;
wire Xd_0__inst_mult_17_28_sumout ;
wire Xd_0__inst_mult_17_29 ;
wire Xd_0__inst_mult_16_263 ;
wire Xd_0__inst_mult_16_264 ;
wire Xd_0__inst_mult_15_258 ;
wire Xd_0__inst_mult_15_259 ;
wire Xd_0__inst_mult_15_28_sumout ;
wire Xd_0__inst_mult_15_29 ;
wire Xd_0__inst_mult_14_253 ;
wire Xd_0__inst_mult_14_254 ;
wire Xd_0__inst_mult_13_253 ;
wire Xd_0__inst_mult_13_254 ;
wire Xd_0__inst_mult_12_253 ;
wire Xd_0__inst_mult_12_254 ;
wire Xd_0__inst_mult_11_253 ;
wire Xd_0__inst_mult_11_254 ;
wire Xd_0__inst_mult_10_253 ;
wire Xd_0__inst_mult_10_254 ;
wire Xd_0__inst_mult_9_253 ;
wire Xd_0__inst_mult_9_254 ;
wire Xd_0__inst_mult_8_253 ;
wire Xd_0__inst_mult_8_254 ;
wire Xd_0__inst_mult_7_253 ;
wire Xd_0__inst_mult_7_254 ;
wire Xd_0__inst_mult_6_253 ;
wire Xd_0__inst_mult_6_254 ;
wire Xd_0__inst_mult_5_253 ;
wire Xd_0__inst_mult_5_254 ;
wire Xd_0__inst_mult_4_239 ;
wire Xd_0__inst_mult_4_240 ;
wire Xd_0__inst_mult_3_234 ;
wire Xd_0__inst_mult_3_235 ;
wire Xd_0__inst_mult_2_229 ;
wire Xd_0__inst_mult_2_230 ;
wire Xd_0__inst_mult_1_234 ;
wire Xd_0__inst_mult_1_235 ;
wire Xd_0__inst_mult_0_234 ;
wire Xd_0__inst_mult_0_235 ;
wire Xd_0__inst_mult_31_234 ;
wire Xd_0__inst_mult_31_33_sumout ;
wire Xd_0__inst_mult_31_34 ;
wire Xd_0__inst_mult_30_249 ;
wire Xd_0__inst_mult_30_250 ;
wire Xd_0__inst_mult_30_33_sumout ;
wire Xd_0__inst_mult_30_34 ;
wire Xd_0__inst_mult_29_234 ;
wire Xd_0__inst_mult_29_33_sumout ;
wire Xd_0__inst_mult_29_34 ;
wire Xd_0__inst_mult_28_239 ;
wire Xd_0__inst_mult_28_240 ;
wire Xd_0__inst_mult_28_33_sumout ;
wire Xd_0__inst_mult_28_34 ;
wire Xd_0__inst_mult_27_234 ;
wire Xd_0__inst_mult_27_33_sumout ;
wire Xd_0__inst_mult_27_34 ;
wire Xd_0__inst_mult_26_249 ;
wire Xd_0__inst_mult_26_250 ;
wire Xd_0__inst_mult_26_33_sumout ;
wire Xd_0__inst_mult_26_34 ;
wire Xd_0__inst_mult_25_244 ;
wire Xd_0__inst_mult_25_33_sumout ;
wire Xd_0__inst_mult_25_34 ;
wire Xd_0__inst_mult_24_244 ;
wire Xd_0__inst_mult_24_245 ;
wire Xd_0__inst_mult_24_33_sumout ;
wire Xd_0__inst_mult_24_34 ;
wire Xd_0__inst_mult_23_254 ;
wire Xd_0__inst_mult_22_254 ;
wire Xd_0__inst_mult_22_255 ;
wire Xd_0__inst_mult_21_254 ;
wire Xd_0__inst_mult_21_33_sumout ;
wire Xd_0__inst_mult_21_34 ;
wire Xd_0__inst_mult_20_268 ;
wire Xd_0__inst_mult_20_269 ;
wire Xd_0__inst_mult_20_33_sumout ;
wire Xd_0__inst_mult_20_34 ;
wire Xd_0__inst_mult_19_268 ;
wire Xd_0__inst_mult_19_33_sumout ;
wire Xd_0__inst_mult_19_34 ;
wire Xd_0__inst_mult_18_268 ;
wire Xd_0__inst_mult_18_269 ;
wire Xd_0__inst_mult_18_33_sumout ;
wire Xd_0__inst_mult_18_34 ;
wire Xd_0__inst_mult_17_268 ;
wire Xd_0__inst_mult_17_33_sumout ;
wire Xd_0__inst_mult_17_34 ;
wire Xd_0__inst_mult_16_268 ;
wire Xd_0__inst_mult_16_269 ;
wire Xd_0__inst_mult_16_33_sumout ;
wire Xd_0__inst_mult_16_34 ;
wire Xd_0__inst_mult_15_263 ;
wire Xd_0__inst_mult_15_33_sumout ;
wire Xd_0__inst_mult_15_34 ;
wire Xd_0__inst_mult_14_258 ;
wire Xd_0__inst_mult_14_259 ;
wire Xd_0__inst_mult_14_33_sumout ;
wire Xd_0__inst_mult_14_34 ;
wire Xd_0__inst_mult_13_258 ;
wire Xd_0__inst_mult_13_33_sumout ;
wire Xd_0__inst_mult_13_34 ;
wire Xd_0__inst_mult_12_258 ;
wire Xd_0__inst_mult_12_259 ;
wire Xd_0__inst_mult_12_33_sumout ;
wire Xd_0__inst_mult_12_34 ;
wire Xd_0__inst_mult_11_258 ;
wire Xd_0__inst_mult_11_33_sumout ;
wire Xd_0__inst_mult_11_34 ;
wire Xd_0__inst_mult_10_258 ;
wire Xd_0__inst_mult_10_259 ;
wire Xd_0__inst_mult_9_258 ;
wire Xd_0__inst_mult_9_33_sumout ;
wire Xd_0__inst_mult_9_34 ;
wire Xd_0__inst_mult_8_258 ;
wire Xd_0__inst_mult_8_259 ;
wire Xd_0__inst_mult_8_33_sumout ;
wire Xd_0__inst_mult_8_34 ;
wire Xd_0__inst_mult_7_258 ;
wire Xd_0__inst_mult_7_33_sumout ;
wire Xd_0__inst_mult_7_34 ;
wire Xd_0__inst_mult_6_258 ;
wire Xd_0__inst_mult_6_259 ;
wire Xd_0__inst_mult_6_33_sumout ;
wire Xd_0__inst_mult_6_34 ;
wire Xd_0__inst_mult_5_258 ;
wire Xd_0__inst_mult_4_244 ;
wire Xd_0__inst_mult_4_245 ;
wire Xd_0__inst_mult_4_33_sumout ;
wire Xd_0__inst_mult_4_34 ;
wire Xd_0__inst_mult_3_239 ;
wire Xd_0__inst_mult_3_33_sumout ;
wire Xd_0__inst_mult_3_34 ;
wire Xd_0__inst_mult_2_234 ;
wire Xd_0__inst_mult_2_235 ;
wire Xd_0__inst_mult_2_33_sumout ;
wire Xd_0__inst_mult_2_34 ;
wire Xd_0__inst_mult_1_239 ;
wire Xd_0__inst_mult_1_33_sumout ;
wire Xd_0__inst_mult_1_34 ;
wire Xd_0__inst_mult_0_239 ;
wire Xd_0__inst_mult_0_240 ;
wire Xd_0__inst_mult_0_33_sumout ;
wire Xd_0__inst_mult_0_34 ;
wire Xd_0__inst_mult_15_268 ;
wire Xd_0__inst_mult_15_269 ;
wire Xd_0__inst_mult_30_254 ;
wire Xd_0__inst_mult_30_255 ;
wire Xd_0__inst_mult_28_244 ;
wire Xd_0__inst_mult_28_245 ;
wire Xd_0__inst_mult_0_244 ;
wire Xd_0__inst_mult_0_245 ;
wire Xd_0__inst_mult_26_254 ;
wire Xd_0__inst_mult_26_255 ;
wire Xd_0__inst_mult_3_244 ;
wire Xd_0__inst_mult_3_245 ;
wire Xd_0__inst_mult_1_244 ;
wire Xd_0__inst_mult_1_245 ;
wire Xd_0__inst_mult_31_239 ;
wire Xd_0__inst_mult_31_240 ;
wire Xd_0__inst_mult_31_245 ;
wire Xd_0__inst_mult_23_259 ;
wire Xd_0__inst_mult_23_260 ;
wire Xd_0__inst_mult_30_259 ;
wire Xd_0__inst_mult_30_260 ;
wire Xd_0__inst_mult_30_265 ;
wire Xd_0__inst_mult_22_259 ;
wire Xd_0__inst_mult_22_260 ;
wire Xd_0__inst_mult_29_239 ;
wire Xd_0__inst_mult_29_240 ;
wire Xd_0__inst_mult_29_245 ;
wire Xd_0__inst_mult_21_259 ;
wire Xd_0__inst_mult_21_260 ;
wire Xd_0__inst_mult_28_249 ;
wire Xd_0__inst_mult_28_250 ;
wire Xd_0__inst_mult_28_255 ;
wire Xd_0__inst_mult_20_273 ;
wire Xd_0__inst_mult_20_274 ;
wire Xd_0__inst_mult_27_239 ;
wire Xd_0__inst_mult_27_240 ;
wire Xd_0__inst_mult_27_245 ;
wire Xd_0__inst_mult_25_249 ;
wire Xd_0__inst_mult_25_250 ;
wire Xd_0__inst_mult_26_259 ;
wire Xd_0__inst_mult_26_260 ;
wire Xd_0__inst_mult_26_265 ;
wire Xd_0__inst_mult_19_273 ;
wire Xd_0__inst_mult_19_274 ;
wire Xd_0__inst_mult_25_254 ;
wire Xd_0__inst_mult_25_255 ;
wire Xd_0__inst_mult_25_260 ;
wire Xd_0__inst_mult_18_273 ;
wire Xd_0__inst_mult_18_274 ;
wire Xd_0__inst_mult_24_249 ;
wire Xd_0__inst_mult_24_250 ;
wire Xd_0__inst_mult_24_255 ;
wire Xd_0__inst_mult_17_273 ;
wire Xd_0__inst_mult_17_274 ;
wire Xd_0__inst_mult_23_264 ;
wire Xd_0__inst_mult_23_265 ;
wire Xd_0__inst_mult_23_270 ;
wire Xd_0__inst_mult_24_259 ;
wire Xd_0__inst_mult_24_260 ;
wire Xd_0__inst_mult_22_264 ;
wire Xd_0__inst_mult_22_265 ;
wire Xd_0__inst_mult_22_270 ;
wire Xd_0__inst_mult_4_249 ;
wire Xd_0__inst_mult_4_250 ;
wire Xd_0__inst_mult_21_264 ;
wire Xd_0__inst_mult_21_265 ;
wire Xd_0__inst_mult_21_270 ;
wire Xd_0__inst_mult_26_269 ;
wire Xd_0__inst_mult_26_270 ;
wire Xd_0__inst_mult_20_278 ;
wire Xd_0__inst_mult_20_279 ;
wire Xd_0__inst_mult_20_284 ;
wire Xd_0__inst_mult_16_273 ;
wire Xd_0__inst_mult_16_274 ;
wire Xd_0__inst_mult_19_278 ;
wire Xd_0__inst_mult_19_279 ;
wire Xd_0__inst_mult_19_284 ;
wire Xd_0__inst_mult_12_263 ;
wire Xd_0__inst_mult_12_264 ;
wire Xd_0__inst_mult_18_278 ;
wire Xd_0__inst_mult_18_279 ;
wire Xd_0__inst_mult_18_284 ;
wire Xd_0__inst_mult_23_274 ;
wire Xd_0__inst_mult_23_275 ;
wire Xd_0__inst_mult_17_278 ;
wire Xd_0__inst_mult_17_279 ;
wire Xd_0__inst_mult_17_284 ;
wire Xd_0__inst_mult_5_263 ;
wire Xd_0__inst_mult_5_264 ;
wire Xd_0__inst_mult_16_278 ;
wire Xd_0__inst_mult_16_279 ;
wire Xd_0__inst_mult_16_284 ;
wire Xd_0__inst_mult_6_263 ;
wire Xd_0__inst_mult_6_264 ;
wire Xd_0__inst_mult_15_273 ;
wire Xd_0__inst_mult_15_274 ;
wire Xd_0__inst_mult_15_279 ;
wire Xd_0__inst_mult_7_263 ;
wire Xd_0__inst_mult_7_264 ;
wire Xd_0__inst_mult_14_263 ;
wire Xd_0__inst_mult_14_264 ;
wire Xd_0__inst_mult_14_269 ;
wire Xd_0__inst_mult_8_263 ;
wire Xd_0__inst_mult_8_264 ;
wire Xd_0__inst_mult_13_263 ;
wire Xd_0__inst_mult_13_264 ;
wire Xd_0__inst_mult_13_269 ;
wire Xd_0__inst_mult_9_263 ;
wire Xd_0__inst_mult_9_264 ;
wire Xd_0__inst_mult_12_268 ;
wire Xd_0__inst_mult_12_269 ;
wire Xd_0__inst_mult_12_274 ;
wire Xd_0__inst_mult_19_288 ;
wire Xd_0__inst_mult_19_289 ;
wire Xd_0__inst_mult_11_263 ;
wire Xd_0__inst_mult_11_264 ;
wire Xd_0__inst_mult_11_269 ;
wire Xd_0__inst_mult_10_263 ;
wire Xd_0__inst_mult_10_264 ;
wire Xd_0__inst_mult_10_268 ;
wire Xd_0__inst_mult_10_269 ;
wire Xd_0__inst_mult_10_274 ;
wire Xd_0__inst_mult_11_273 ;
wire Xd_0__inst_mult_11_274 ;
wire Xd_0__inst_mult_9_268 ;
wire Xd_0__inst_mult_9_269 ;
wire Xd_0__inst_mult_9_274 ;
wire Xd_0__inst_mult_13_273 ;
wire Xd_0__inst_mult_13_274 ;
wire Xd_0__inst_mult_8_268 ;
wire Xd_0__inst_mult_8_269 ;
wire Xd_0__inst_mult_8_274 ;
wire Xd_0__inst_mult_14_273 ;
wire Xd_0__inst_mult_14_274 ;
wire Xd_0__inst_mult_7_268 ;
wire Xd_0__inst_mult_7_269 ;
wire Xd_0__inst_mult_7_274 ;
wire Xd_0__inst_mult_15_283 ;
wire Xd_0__inst_mult_15_284 ;
wire Xd_0__inst_mult_6_268 ;
wire Xd_0__inst_mult_6_269 ;
wire Xd_0__inst_mult_6_274 ;
wire Xd_0__inst_mult_16_288 ;
wire Xd_0__inst_mult_16_289 ;
wire Xd_0__inst_mult_5_268 ;
wire Xd_0__inst_mult_5_269 ;
wire Xd_0__inst_mult_5_274 ;
wire Xd_0__inst_mult_17_288 ;
wire Xd_0__inst_mult_17_289 ;
wire Xd_0__inst_mult_4_254 ;
wire Xd_0__inst_mult_4_255 ;
wire Xd_0__inst_mult_4_260 ;
wire Xd_0__inst_mult_18_288 ;
wire Xd_0__inst_mult_18_289 ;
wire Xd_0__inst_mult_3_249 ;
wire Xd_0__inst_mult_3_250 ;
wire Xd_0__inst_mult_3_255 ;
wire Xd_0__inst_mult_30_269 ;
wire Xd_0__inst_mult_30_270 ;
wire Xd_0__inst_mult_2_239 ;
wire Xd_0__inst_mult_2_240 ;
wire Xd_0__inst_mult_2_245 ;
wire Xd_0__inst_mult_20_288 ;
wire Xd_0__inst_mult_20_289 ;
wire Xd_0__inst_mult_1_249 ;
wire Xd_0__inst_mult_1_250 ;
wire Xd_0__inst_mult_1_255 ;
wire Xd_0__inst_mult_21_274 ;
wire Xd_0__inst_mult_21_275 ;
wire Xd_0__inst_mult_0_249 ;
wire Xd_0__inst_mult_0_250 ;
wire Xd_0__inst_mult_0_255 ;
wire Xd_0__inst_mult_22_274 ;
wire Xd_0__inst_mult_22_275 ;
wire Xd_0__inst_mult_31_249 ;
wire Xd_0__inst_mult_31_250 ;
wire Xd_0__inst_mult_30_274 ;
wire Xd_0__inst_mult_30_275 ;
wire Xd_0__inst_mult_29_249 ;
wire Xd_0__inst_mult_29_250 ;
wire Xd_0__inst_mult_31_254 ;
wire Xd_0__inst_mult_31_255 ;
wire Xd_0__inst_mult_28_259 ;
wire Xd_0__inst_mult_28_260 ;
wire Xd_0__inst_mult_27_249 ;
wire Xd_0__inst_mult_27_250 ;
wire Xd_0__inst_mult_28_264 ;
wire Xd_0__inst_mult_28_265 ;
wire Xd_0__inst_mult_26_274 ;
wire Xd_0__inst_mult_26_275 ;
wire Xd_0__inst_mult_25_264 ;
wire Xd_0__inst_mult_25_265 ;
wire Xd_0__inst_mult_24_264 ;
wire Xd_0__inst_mult_24_265 ;
wire Xd_0__inst_mult_23_279 ;
wire Xd_0__inst_mult_23_280 ;
wire Xd_0__inst_mult_22_279 ;
wire Xd_0__inst_mult_22_280 ;
wire Xd_0__inst_mult_21_279 ;
wire Xd_0__inst_mult_21_280 ;
wire Xd_0__inst_mult_20_293 ;
wire Xd_0__inst_mult_20_294 ;
wire Xd_0__inst_mult_19_293 ;
wire Xd_0__inst_mult_19_294 ;
wire Xd_0__inst_mult_18_293 ;
wire Xd_0__inst_mult_18_294 ;
wire Xd_0__inst_mult_17_293 ;
wire Xd_0__inst_mult_17_294 ;
wire Xd_0__inst_mult_16_293 ;
wire Xd_0__inst_mult_16_294 ;
wire Xd_0__inst_mult_15_288 ;
wire Xd_0__inst_mult_15_289 ;
wire Xd_0__inst_mult_14_278 ;
wire Xd_0__inst_mult_14_279 ;
wire Xd_0__inst_mult_13_278 ;
wire Xd_0__inst_mult_13_279 ;
wire Xd_0__inst_mult_13_283 ;
wire Xd_0__inst_mult_13_284 ;
wire Xd_0__inst_mult_12_278 ;
wire Xd_0__inst_mult_12_279 ;
wire Xd_0__inst_mult_11_278 ;
wire Xd_0__inst_mult_11_279 ;
wire Xd_0__inst_mult_11_283 ;
wire Xd_0__inst_mult_11_284 ;
wire Xd_0__inst_mult_10_278 ;
wire Xd_0__inst_mult_10_279 ;
wire Xd_0__inst_mult_9_278 ;
wire Xd_0__inst_mult_9_279 ;
wire Xd_0__inst_mult_10_283 ;
wire Xd_0__inst_mult_10_284 ;
wire Xd_0__inst_mult_8_278 ;
wire Xd_0__inst_mult_8_279 ;
wire Xd_0__inst_mult_7_278 ;
wire Xd_0__inst_mult_7_279 ;
wire Xd_0__inst_mult_8_283 ;
wire Xd_0__inst_mult_8_284 ;
wire Xd_0__inst_mult_6_278 ;
wire Xd_0__inst_mult_6_279 ;
wire Xd_0__inst_mult_5_278 ;
wire Xd_0__inst_mult_5_279 ;
wire Xd_0__inst_mult_6_283 ;
wire Xd_0__inst_mult_6_284 ;
wire Xd_0__inst_mult_4_264 ;
wire Xd_0__inst_mult_4_265 ;
wire Xd_0__inst_mult_3_259 ;
wire Xd_0__inst_mult_3_260 ;
wire Xd_0__inst_mult_4_269 ;
wire Xd_0__inst_mult_4_270 ;
wire Xd_0__inst_mult_2_249 ;
wire Xd_0__inst_mult_2_250 ;
wire Xd_0__inst_mult_1_259 ;
wire Xd_0__inst_mult_1_260 ;
wire Xd_0__inst_mult_2_254 ;
wire Xd_0__inst_mult_2_255 ;
wire Xd_0__inst_mult_0_259 ;
wire Xd_0__inst_mult_0_260 ;
wire Xd_0__inst_mult_31_259 ;
wire Xd_0__inst_mult_31_260 ;
wire Xd_0__inst_mult_30_279 ;
wire Xd_0__inst_mult_30_280 ;
wire Xd_0__inst_mult_29_254 ;
wire Xd_0__inst_mult_29_255 ;
wire Xd_0__inst_mult_28_269 ;
wire Xd_0__inst_mult_28_270 ;
wire Xd_0__inst_mult_27_254 ;
wire Xd_0__inst_mult_27_255 ;
wire Xd_0__inst_mult_26_279 ;
wire Xd_0__inst_mult_26_280 ;
wire Xd_0__inst_mult_25_269 ;
wire Xd_0__inst_mult_25_270 ;
wire Xd_0__inst_mult_24_269 ;
wire Xd_0__inst_mult_24_270 ;
wire Xd_0__inst_mult_23_284 ;
wire Xd_0__inst_mult_23_285 ;
wire Xd_0__inst_mult_22_284 ;
wire Xd_0__inst_mult_22_285 ;
wire Xd_0__inst_mult_21_284 ;
wire Xd_0__inst_mult_21_285 ;
wire Xd_0__inst_mult_20_298 ;
wire Xd_0__inst_mult_20_299 ;
wire Xd_0__inst_mult_19_298 ;
wire Xd_0__inst_mult_19_299 ;
wire Xd_0__inst_mult_18_298 ;
wire Xd_0__inst_mult_18_299 ;
wire Xd_0__inst_mult_17_298 ;
wire Xd_0__inst_mult_17_299 ;
wire Xd_0__inst_mult_16_298 ;
wire Xd_0__inst_mult_16_299 ;
wire Xd_0__inst_mult_15_293 ;
wire Xd_0__inst_mult_15_294 ;
wire Xd_0__inst_mult_14_283 ;
wire Xd_0__inst_mult_14_284 ;
wire Xd_0__inst_mult_13_288 ;
wire Xd_0__inst_mult_13_289 ;
wire Xd_0__inst_mult_12_283 ;
wire Xd_0__inst_mult_12_284 ;
wire Xd_0__inst_mult_11_288 ;
wire Xd_0__inst_mult_11_289 ;
wire Xd_0__inst_mult_10_288 ;
wire Xd_0__inst_mult_10_289 ;
wire Xd_0__inst_mult_9_283 ;
wire Xd_0__inst_mult_9_284 ;
wire Xd_0__inst_mult_8_288 ;
wire Xd_0__inst_mult_8_289 ;
wire Xd_0__inst_mult_7_283 ;
wire Xd_0__inst_mult_7_284 ;
wire Xd_0__inst_mult_6_288 ;
wire Xd_0__inst_mult_6_289 ;
wire Xd_0__inst_mult_5_283 ;
wire Xd_0__inst_mult_5_284 ;
wire Xd_0__inst_mult_4_274 ;
wire Xd_0__inst_mult_4_275 ;
wire Xd_0__inst_mult_3_264 ;
wire Xd_0__inst_mult_3_265 ;
wire Xd_0__inst_mult_2_259 ;
wire Xd_0__inst_mult_2_260 ;
wire Xd_0__inst_mult_1_264 ;
wire Xd_0__inst_mult_1_265 ;
wire Xd_0__inst_mult_0_264 ;
wire Xd_0__inst_mult_0_265 ;
wire Xd_0__inst_mult_31_264 ;
wire Xd_0__inst_mult_31_265 ;
wire Xd_0__inst_mult_31_269 ;
wire Xd_0__inst_mult_31_270 ;
wire Xd_0__inst_mult_31_274 ;
wire Xd_0__inst_mult_31_275 ;
wire Xd_0__inst_mult_31_280 ;
wire Xd_0__inst_mult_30_284 ;
wire Xd_0__inst_mult_30_285 ;
wire Xd_0__inst_mult_30_289 ;
wire Xd_0__inst_mult_30_290 ;
wire Xd_0__inst_mult_30_294 ;
wire Xd_0__inst_mult_30_295 ;
wire Xd_0__inst_mult_30_300 ;
wire Xd_0__inst_mult_29_259 ;
wire Xd_0__inst_mult_29_260 ;
wire Xd_0__inst_mult_29_264 ;
wire Xd_0__inst_mult_29_265 ;
wire Xd_0__inst_mult_29_269 ;
wire Xd_0__inst_mult_29_270 ;
wire Xd_0__inst_mult_29_275 ;
wire Xd_0__inst_mult_28_274 ;
wire Xd_0__inst_mult_28_275 ;
wire Xd_0__inst_mult_28_279 ;
wire Xd_0__inst_mult_28_280 ;
wire Xd_0__inst_mult_28_284 ;
wire Xd_0__inst_mult_28_285 ;
wire Xd_0__inst_mult_28_290 ;
wire Xd_0__inst_mult_27_259 ;
wire Xd_0__inst_mult_27_260 ;
wire Xd_0__inst_mult_27_264 ;
wire Xd_0__inst_mult_27_265 ;
wire Xd_0__inst_mult_27_269 ;
wire Xd_0__inst_mult_27_270 ;
wire Xd_0__inst_mult_27_275 ;
wire Xd_0__inst_mult_26_284 ;
wire Xd_0__inst_mult_26_285 ;
wire Xd_0__inst_mult_26_289 ;
wire Xd_0__inst_mult_26_290 ;
wire Xd_0__inst_mult_26_294 ;
wire Xd_0__inst_mult_26_295 ;
wire Xd_0__inst_mult_26_300 ;
wire Xd_0__inst_mult_25_274 ;
wire Xd_0__inst_mult_25_275 ;
wire Xd_0__inst_mult_25_279 ;
wire Xd_0__inst_mult_25_280 ;
wire Xd_0__inst_mult_25_284 ;
wire Xd_0__inst_mult_25_285 ;
wire Xd_0__inst_mult_25_290 ;
wire Xd_0__inst_mult_24_274 ;
wire Xd_0__inst_mult_24_275 ;
wire Xd_0__inst_mult_24_279 ;
wire Xd_0__inst_mult_24_280 ;
wire Xd_0__inst_mult_24_284 ;
wire Xd_0__inst_mult_24_285 ;
wire Xd_0__inst_mult_24_290 ;
wire Xd_0__inst_mult_23_289 ;
wire Xd_0__inst_mult_23_290 ;
wire Xd_0__inst_mult_23_294 ;
wire Xd_0__inst_mult_23_295 ;
wire Xd_0__inst_mult_23_300 ;
wire Xd_0__inst_mult_22_289 ;
wire Xd_0__inst_mult_22_290 ;
wire Xd_0__inst_mult_22_294 ;
wire Xd_0__inst_mult_22_295 ;
wire Xd_0__inst_mult_22_300 ;
wire Xd_0__inst_mult_21_289 ;
wire Xd_0__inst_mult_21_290 ;
wire Xd_0__inst_mult_21_294 ;
wire Xd_0__inst_mult_21_295 ;
wire Xd_0__inst_mult_21_300 ;
wire Xd_0__inst_mult_20_303 ;
wire Xd_0__inst_mult_20_304 ;
wire Xd_0__inst_mult_20_309 ;
wire Xd_0__inst_mult_19_303 ;
wire Xd_0__inst_mult_19_304 ;
wire Xd_0__inst_mult_19_309 ;
wire Xd_0__inst_mult_18_303 ;
wire Xd_0__inst_mult_18_304 ;
wire Xd_0__inst_mult_18_309 ;
wire Xd_0__inst_mult_17_303 ;
wire Xd_0__inst_mult_17_304 ;
wire Xd_0__inst_mult_17_309 ;
wire Xd_0__inst_mult_16_303 ;
wire Xd_0__inst_mult_16_304 ;
wire Xd_0__inst_mult_16_309 ;
wire Xd_0__inst_mult_15_298 ;
wire Xd_0__inst_mult_15_299 ;
wire Xd_0__inst_mult_15_304 ;
wire Xd_0__inst_mult_14_288 ;
wire Xd_0__inst_mult_14_289 ;
wire Xd_0__inst_mult_14_294 ;
wire Xd_0__inst_mult_13_293 ;
wire Xd_0__inst_mult_13_294 ;
wire Xd_0__inst_mult_13_299 ;
wire Xd_0__inst_mult_12_288 ;
wire Xd_0__inst_mult_12_289 ;
wire Xd_0__inst_mult_12_294 ;
wire Xd_0__inst_mult_11_293 ;
wire Xd_0__inst_mult_11_294 ;
wire Xd_0__inst_mult_11_299 ;
wire Xd_0__inst_mult_10_293 ;
wire Xd_0__inst_mult_10_294 ;
wire Xd_0__inst_mult_10_299 ;
wire Xd_0__inst_mult_9_288 ;
wire Xd_0__inst_mult_9_289 ;
wire Xd_0__inst_mult_9_294 ;
wire Xd_0__inst_mult_8_293 ;
wire Xd_0__inst_mult_8_294 ;
wire Xd_0__inst_mult_8_299 ;
wire Xd_0__inst_mult_7_288 ;
wire Xd_0__inst_mult_7_289 ;
wire Xd_0__inst_mult_7_294 ;
wire Xd_0__inst_mult_6_293 ;
wire Xd_0__inst_mult_6_294 ;
wire Xd_0__inst_mult_6_299 ;
wire Xd_0__inst_mult_5_288 ;
wire Xd_0__inst_mult_5_289 ;
wire Xd_0__inst_mult_5_294 ;
wire Xd_0__inst_mult_4_279 ;
wire Xd_0__inst_mult_4_280 ;
wire Xd_0__inst_mult_4_284 ;
wire Xd_0__inst_mult_4_285 ;
wire Xd_0__inst_mult_4_290 ;
wire Xd_0__inst_mult_3_269 ;
wire Xd_0__inst_mult_3_270 ;
wire Xd_0__inst_mult_3_274 ;
wire Xd_0__inst_mult_3_275 ;
wire Xd_0__inst_mult_3_279 ;
wire Xd_0__inst_mult_3_280 ;
wire Xd_0__inst_mult_3_285 ;
wire Xd_0__inst_mult_2_264 ;
wire Xd_0__inst_mult_2_265 ;
wire Xd_0__inst_mult_2_269 ;
wire Xd_0__inst_mult_2_270 ;
wire Xd_0__inst_mult_2_274 ;
wire Xd_0__inst_mult_2_275 ;
wire Xd_0__inst_mult_2_280 ;
wire Xd_0__inst_mult_1_269 ;
wire Xd_0__inst_mult_1_270 ;
wire Xd_0__inst_mult_1_274 ;
wire Xd_0__inst_mult_1_275 ;
wire Xd_0__inst_mult_1_279 ;
wire Xd_0__inst_mult_1_280 ;
wire Xd_0__inst_mult_1_285 ;
wire Xd_0__inst_mult_0_269 ;
wire Xd_0__inst_mult_0_270 ;
wire Xd_0__inst_mult_0_274 ;
wire Xd_0__inst_mult_0_275 ;
wire Xd_0__inst_mult_0_279 ;
wire Xd_0__inst_mult_0_280 ;
wire Xd_0__inst_mult_0_285 ;
wire Xd_0__inst_mult_31_284 ;
wire Xd_0__inst_mult_31_285 ;
wire Xd_0__inst_mult_31_289 ;
wire Xd_0__inst_mult_31_290 ;
wire Xd_0__inst_mult_31_294 ;
wire Xd_0__inst_mult_31_295 ;
wire Xd_0__inst_mult_30_304 ;
wire Xd_0__inst_mult_30_305 ;
wire Xd_0__inst_mult_30_309 ;
wire Xd_0__inst_mult_30_310 ;
wire Xd_0__inst_mult_29_279 ;
wire Xd_0__inst_mult_29_280 ;
wire Xd_0__inst_mult_29_284 ;
wire Xd_0__inst_mult_29_285 ;
wire Xd_0__inst_mult_29_289 ;
wire Xd_0__inst_mult_29_290 ;
wire Xd_0__inst_mult_28_294 ;
wire Xd_0__inst_mult_28_295 ;
wire Xd_0__inst_mult_28_299 ;
wire Xd_0__inst_mult_28_300 ;
wire Xd_0__inst_mult_27_279 ;
wire Xd_0__inst_mult_27_280 ;
wire Xd_0__inst_mult_27_284 ;
wire Xd_0__inst_mult_27_285 ;
wire Xd_0__inst_mult_27_289 ;
wire Xd_0__inst_mult_27_290 ;
wire Xd_0__inst_mult_26_304 ;
wire Xd_0__inst_mult_26_305 ;
wire Xd_0__inst_mult_26_309 ;
wire Xd_0__inst_mult_26_310 ;
wire Xd_0__inst_mult_25_294 ;
wire Xd_0__inst_mult_25_295 ;
wire Xd_0__inst_mult_25_299 ;
wire Xd_0__inst_mult_25_300 ;
wire Xd_0__inst_mult_25_304 ;
wire Xd_0__inst_mult_25_305 ;
wire Xd_0__inst_mult_24_294 ;
wire Xd_0__inst_mult_24_295 ;
wire Xd_0__inst_mult_24_299 ;
wire Xd_0__inst_mult_24_300 ;
wire Xd_0__inst_mult_24_304 ;
wire Xd_0__inst_mult_24_305 ;
wire Xd_0__inst_mult_23_304 ;
wire Xd_0__inst_mult_23_305 ;
wire Xd_0__inst_mult_23_309 ;
wire Xd_0__inst_mult_23_310 ;
wire Xd_0__inst_mult_22_304 ;
wire Xd_0__inst_mult_22_305 ;
wire Xd_0__inst_mult_22_309 ;
wire Xd_0__inst_mult_22_310 ;
wire Xd_0__inst_mult_21_304 ;
wire Xd_0__inst_mult_21_305 ;
wire Xd_0__inst_mult_21_309 ;
wire Xd_0__inst_mult_21_310 ;
wire Xd_0__inst_mult_20_313 ;
wire Xd_0__inst_mult_20_314 ;
wire Xd_0__inst_mult_19_313 ;
wire Xd_0__inst_mult_19_314 ;
wire Xd_0__inst_mult_18_313 ;
wire Xd_0__inst_mult_18_314 ;
wire Xd_0__inst_mult_17_313 ;
wire Xd_0__inst_mult_17_314 ;
wire Xd_0__inst_mult_16_313 ;
wire Xd_0__inst_mult_16_314 ;
wire Xd_0__inst_mult_15_308 ;
wire Xd_0__inst_mult_15_309 ;
wire Xd_0__inst_mult_14_298 ;
wire Xd_0__inst_mult_14_299 ;
wire Xd_0__inst_mult_13_303 ;
wire Xd_0__inst_mult_13_304 ;
wire Xd_0__inst_mult_12_298 ;
wire Xd_0__inst_mult_12_299 ;
wire Xd_0__inst_mult_11_303 ;
wire Xd_0__inst_mult_11_304 ;
wire Xd_0__inst_mult_10_303 ;
wire Xd_0__inst_mult_10_304 ;
wire Xd_0__inst_mult_9_298 ;
wire Xd_0__inst_mult_9_299 ;
wire Xd_0__inst_mult_8_303 ;
wire Xd_0__inst_mult_8_304 ;
wire Xd_0__inst_mult_7_298 ;
wire Xd_0__inst_mult_7_299 ;
wire Xd_0__inst_mult_6_303 ;
wire Xd_0__inst_mult_6_304 ;
wire Xd_0__inst_mult_5_298 ;
wire Xd_0__inst_mult_5_299 ;
wire Xd_0__inst_mult_4_294 ;
wire Xd_0__inst_mult_4_295 ;
wire Xd_0__inst_mult_4_299 ;
wire Xd_0__inst_mult_4_300 ;
wire Xd_0__inst_mult_3_289 ;
wire Xd_0__inst_mult_3_290 ;
wire Xd_0__inst_mult_3_294 ;
wire Xd_0__inst_mult_3_295 ;
wire Xd_0__inst_mult_2_284 ;
wire Xd_0__inst_mult_2_285 ;
wire Xd_0__inst_mult_2_289 ;
wire Xd_0__inst_mult_2_290 ;
wire Xd_0__inst_mult_2_294 ;
wire Xd_0__inst_mult_2_295 ;
wire Xd_0__inst_mult_1_289 ;
wire Xd_0__inst_mult_1_290 ;
wire Xd_0__inst_mult_1_294 ;
wire Xd_0__inst_mult_1_295 ;
wire Xd_0__inst_mult_0_289 ;
wire Xd_0__inst_mult_0_290 ;
wire Xd_0__inst_mult_0_294 ;
wire Xd_0__inst_mult_0_295 ;
wire Xd_0__inst_mult_0_299 ;
wire Xd_0__inst_mult_0_300 ;
wire Xd_0__inst_mult_31_299 ;
wire Xd_0__inst_mult_31_304 ;
wire Xd_0__inst_mult_31_305 ;
wire Xd_0__inst_mult_31_309 ;
wire Xd_0__inst_mult_31_310 ;
wire Xd_0__inst_mult_30_314 ;
wire Xd_0__inst_mult_30_315 ;
wire Xd_0__inst_mult_30_319 ;
wire Xd_0__inst_mult_30_320 ;
wire Xd_0__inst_mult_29_294 ;
wire Xd_0__inst_mult_29_299 ;
wire Xd_0__inst_mult_29_300 ;
wire Xd_0__inst_mult_29_304 ;
wire Xd_0__inst_mult_29_305 ;
wire Xd_0__inst_mult_28_304 ;
wire Xd_0__inst_mult_28_305 ;
wire Xd_0__inst_mult_28_309 ;
wire Xd_0__inst_mult_28_310 ;
wire Xd_0__inst_mult_27_294 ;
wire Xd_0__inst_mult_27_299 ;
wire Xd_0__inst_mult_27_300 ;
wire Xd_0__inst_mult_27_304 ;
wire Xd_0__inst_mult_27_305 ;
wire Xd_0__inst_mult_26_314 ;
wire Xd_0__inst_mult_26_315 ;
wire Xd_0__inst_mult_26_319 ;
wire Xd_0__inst_mult_26_320 ;
wire Xd_0__inst_mult_25_309 ;
wire Xd_0__inst_mult_25_314 ;
wire Xd_0__inst_mult_25_315 ;
wire Xd_0__inst_mult_25_319 ;
wire Xd_0__inst_mult_25_320 ;
wire Xd_0__inst_mult_24_309 ;
wire Xd_0__inst_mult_24_314 ;
wire Xd_0__inst_mult_24_315 ;
wire Xd_0__inst_mult_24_319 ;
wire Xd_0__inst_mult_24_320 ;
wire Xd_0__inst_mult_23_314 ;
wire Xd_0__inst_mult_23_315 ;
wire Xd_0__inst_mult_23_319 ;
wire Xd_0__inst_mult_23_320 ;
wire Xd_0__inst_mult_22_314 ;
wire Xd_0__inst_mult_22_315 ;
wire Xd_0__inst_mult_22_319 ;
wire Xd_0__inst_mult_22_320 ;
wire Xd_0__inst_mult_21_314 ;
wire Xd_0__inst_mult_21_315 ;
wire Xd_0__inst_mult_21_319 ;
wire Xd_0__inst_mult_21_320 ;
wire Xd_0__inst_mult_20_318 ;
wire Xd_0__inst_mult_20_319 ;
wire Xd_0__inst_mult_19_318 ;
wire Xd_0__inst_mult_19_319 ;
wire Xd_0__inst_mult_18_318 ;
wire Xd_0__inst_mult_18_319 ;
wire Xd_0__inst_mult_17_318 ;
wire Xd_0__inst_mult_17_319 ;
wire Xd_0__inst_mult_16_318 ;
wire Xd_0__inst_mult_16_319 ;
wire Xd_0__inst_mult_15_313 ;
wire Xd_0__inst_mult_15_314 ;
wire Xd_0__inst_mult_14_303 ;
wire Xd_0__inst_mult_14_304 ;
wire Xd_0__inst_mult_13_308 ;
wire Xd_0__inst_mult_13_309 ;
wire Xd_0__inst_mult_12_303 ;
wire Xd_0__inst_mult_12_304 ;
wire Xd_0__inst_mult_11_308 ;
wire Xd_0__inst_mult_11_309 ;
wire Xd_0__inst_mult_10_308 ;
wire Xd_0__inst_mult_10_309 ;
wire Xd_0__inst_mult_9_303 ;
wire Xd_0__inst_mult_9_304 ;
wire Xd_0__inst_mult_8_308 ;
wire Xd_0__inst_mult_8_309 ;
wire Xd_0__inst_mult_7_303 ;
wire Xd_0__inst_mult_7_304 ;
wire Xd_0__inst_mult_6_308 ;
wire Xd_0__inst_mult_6_309 ;
wire Xd_0__inst_mult_5_303 ;
wire Xd_0__inst_mult_5_304 ;
wire Xd_0__inst_mult_4_304 ;
wire Xd_0__inst_mult_4_305 ;
wire Xd_0__inst_mult_4_309 ;
wire Xd_0__inst_mult_4_310 ;
wire Xd_0__inst_mult_3_299 ;
wire Xd_0__inst_mult_3_300 ;
wire Xd_0__inst_mult_3_304 ;
wire Xd_0__inst_mult_3_305 ;
wire Xd_0__inst_mult_2_299 ;
wire Xd_0__inst_mult_2_304 ;
wire Xd_0__inst_mult_2_305 ;
wire Xd_0__inst_mult_2_309 ;
wire Xd_0__inst_mult_2_310 ;
wire Xd_0__inst_mult_1_299 ;
wire Xd_0__inst_mult_1_300 ;
wire Xd_0__inst_mult_1_304 ;
wire Xd_0__inst_mult_1_305 ;
wire Xd_0__inst_mult_0_304 ;
wire Xd_0__inst_mult_0_309 ;
wire Xd_0__inst_mult_0_310 ;
wire Xd_0__inst_mult_0_314 ;
wire Xd_0__inst_mult_0_315 ;
wire Xd_0__inst_mult_31_314 ;
wire Xd_0__inst_mult_31_315 ;
wire Xd_0__inst_mult_31_319 ;
wire Xd_0__inst_mult_31_320 ;
wire Xd_0__inst_mult_30_324 ;
wire Xd_0__inst_mult_30_325 ;
wire Xd_0__inst_mult_29_309 ;
wire Xd_0__inst_mult_29_310 ;
wire Xd_0__inst_mult_29_314 ;
wire Xd_0__inst_mult_29_315 ;
wire Xd_0__inst_mult_28_314 ;
wire Xd_0__inst_mult_28_315 ;
wire Xd_0__inst_mult_28_319 ;
wire Xd_0__inst_mult_28_320 ;
wire Xd_0__inst_mult_27_309 ;
wire Xd_0__inst_mult_27_310 ;
wire Xd_0__inst_mult_27_314 ;
wire Xd_0__inst_mult_27_315 ;
wire Xd_0__inst_mult_26_324 ;
wire Xd_0__inst_mult_26_325 ;
wire Xd_0__inst_mult_25_324 ;
wire Xd_0__inst_mult_25_325 ;
wire Xd_0__inst_mult_24_324 ;
wire Xd_0__inst_mult_24_325 ;
wire Xd_0__inst_mult_23_324 ;
wire Xd_0__inst_mult_23_325 ;
wire Xd_0__inst_mult_22_324 ;
wire Xd_0__inst_mult_22_325 ;
wire Xd_0__inst_mult_21_324 ;
wire Xd_0__inst_mult_21_325 ;
wire Xd_0__inst_mult_15_318 ;
wire Xd_0__inst_mult_15_319 ;
wire Xd_0__inst_mult_14_308 ;
wire Xd_0__inst_mult_14_309 ;
wire Xd_0__inst_mult_13_313 ;
wire Xd_0__inst_mult_13_314 ;
wire Xd_0__inst_mult_12_308 ;
wire Xd_0__inst_mult_12_309 ;
wire Xd_0__inst_mult_11_313 ;
wire Xd_0__inst_mult_11_314 ;
wire Xd_0__inst_mult_10_313 ;
wire Xd_0__inst_mult_10_314 ;
wire Xd_0__inst_mult_9_308 ;
wire Xd_0__inst_mult_9_309 ;
wire Xd_0__inst_mult_8_313 ;
wire Xd_0__inst_mult_8_314 ;
wire Xd_0__inst_mult_7_308 ;
wire Xd_0__inst_mult_7_309 ;
wire Xd_0__inst_mult_6_313 ;
wire Xd_0__inst_mult_6_314 ;
wire Xd_0__inst_mult_5_308 ;
wire Xd_0__inst_mult_5_309 ;
wire Xd_0__inst_mult_4_314 ;
wire Xd_0__inst_mult_4_315 ;
wire Xd_0__inst_mult_4_319 ;
wire Xd_0__inst_mult_4_320 ;
wire Xd_0__inst_mult_3_309 ;
wire Xd_0__inst_mult_3_310 ;
wire Xd_0__inst_mult_3_314 ;
wire Xd_0__inst_mult_3_315 ;
wire Xd_0__inst_mult_2_314 ;
wire Xd_0__inst_mult_2_315 ;
wire Xd_0__inst_mult_2_319 ;
wire Xd_0__inst_mult_2_320 ;
wire Xd_0__inst_mult_1_309 ;
wire Xd_0__inst_mult_1_310 ;
wire Xd_0__inst_mult_1_314 ;
wire Xd_0__inst_mult_1_315 ;
wire Xd_0__inst_mult_0_319 ;
wire Xd_0__inst_mult_0_320 ;
wire Xd_0__inst_mult_0_324 ;
wire Xd_0__inst_mult_0_325 ;
wire Xd_0__inst_mult_31_324 ;
wire Xd_0__inst_mult_31_325 ;
wire Xd_0__inst_mult_29_319 ;
wire Xd_0__inst_mult_29_320 ;
wire Xd_0__inst_mult_28_324 ;
wire Xd_0__inst_mult_28_325 ;
wire Xd_0__inst_mult_27_319 ;
wire Xd_0__inst_mult_27_320 ;
wire Xd_0__inst_mult_14_313 ;
wire Xd_0__inst_mult_14_314 ;
wire Xd_0__inst_mult_13_318 ;
wire Xd_0__inst_mult_13_319 ;
wire Xd_0__inst_mult_12_313 ;
wire Xd_0__inst_mult_12_314 ;
wire Xd_0__inst_mult_11_318 ;
wire Xd_0__inst_mult_11_319 ;
wire Xd_0__inst_mult_10_318 ;
wire Xd_0__inst_mult_10_319 ;
wire Xd_0__inst_mult_9_313 ;
wire Xd_0__inst_mult_9_314 ;
wire Xd_0__inst_mult_8_318 ;
wire Xd_0__inst_mult_8_319 ;
wire Xd_0__inst_mult_7_313 ;
wire Xd_0__inst_mult_7_314 ;
wire Xd_0__inst_mult_6_318 ;
wire Xd_0__inst_mult_6_319 ;
wire Xd_0__inst_mult_5_313 ;
wire Xd_0__inst_mult_5_314 ;
wire Xd_0__inst_mult_4_324 ;
wire Xd_0__inst_mult_4_325 ;
wire Xd_0__inst_mult_3_319 ;
wire Xd_0__inst_mult_3_320 ;
wire Xd_0__inst_mult_2_324 ;
wire Xd_0__inst_mult_2_325 ;
wire Xd_0__inst_mult_1_319 ;
wire Xd_0__inst_mult_1_320 ;
wire Xd_0__inst_mult_29_324 ;
wire Xd_0__inst_mult_27_324 ;
wire Xd_0__inst_mult_14_318 ;
wire Xd_0__inst_mult_12_318 ;
wire Xd_0__inst_mult_9_318 ;
wire Xd_0__inst_mult_7_318 ;
wire Xd_0__inst_mult_5_318 ;
wire Xd_0__inst_mult_3_324 ;
wire Xd_0__inst_mult_1_324 ;
wire Xd_0__inst_inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_inst_first_level_0__17__q ;
wire Xd_0__inst_inst_inst_first_level_1__18__q ;
wire Xd_0__inst_inst_inst_first_level_0__18__q ;
wire Xd_0__inst_inst_first_level_3__0__q ;
wire Xd_0__inst_inst_first_level_2__0__q ;
wire Xd_0__inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_first_level_3__1__q ;
wire Xd_0__inst_inst_first_level_2__1__q ;
wire Xd_0__inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_first_level_3__2__q ;
wire Xd_0__inst_inst_first_level_2__2__q ;
wire Xd_0__inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_first_level_3__3__q ;
wire Xd_0__inst_inst_first_level_2__3__q ;
wire Xd_0__inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_first_level_3__4__q ;
wire Xd_0__inst_inst_first_level_2__4__q ;
wire Xd_0__inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_first_level_3__5__q ;
wire Xd_0__inst_inst_first_level_2__5__q ;
wire Xd_0__inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_first_level_3__6__q ;
wire Xd_0__inst_inst_first_level_2__6__q ;
wire Xd_0__inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_first_level_3__7__q ;
wire Xd_0__inst_inst_first_level_2__7__q ;
wire Xd_0__inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_first_level_3__8__q ;
wire Xd_0__inst_inst_first_level_2__8__q ;
wire Xd_0__inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_first_level_3__9__q ;
wire Xd_0__inst_inst_first_level_2__9__q ;
wire Xd_0__inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_first_level_3__10__q ;
wire Xd_0__inst_inst_first_level_2__10__q ;
wire Xd_0__inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_first_level_3__11__q ;
wire Xd_0__inst_inst_first_level_2__11__q ;
wire Xd_0__inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_first_level_3__12__q ;
wire Xd_0__inst_inst_first_level_2__12__q ;
wire Xd_0__inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_first_level_3__13__q ;
wire Xd_0__inst_inst_first_level_2__13__q ;
wire Xd_0__inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_first_level_3__14__q ;
wire Xd_0__inst_inst_first_level_2__14__q ;
wire Xd_0__inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_first_level_3__15__q ;
wire Xd_0__inst_inst_first_level_2__15__q ;
wire Xd_0__inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_first_level_3__16__q ;
wire Xd_0__inst_inst_first_level_2__16__q ;
wire Xd_0__inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_first_level_3__17__q ;
wire Xd_0__inst_inst_first_level_2__17__q ;
wire Xd_0__inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_first_level_0__17__q ;
wire Xd_0__inst_r_sum2_7__0__q ;
wire Xd_0__inst_r_sum2_6__0__q ;
wire Xd_0__inst_r_sum2_5__0__q ;
wire Xd_0__inst_r_sum2_4__0__q ;
wire Xd_0__inst_r_sum2_3__0__q ;
wire Xd_0__inst_r_sum2_2__0__q ;
wire Xd_0__inst_r_sum2_1__0__q ;
wire Xd_0__inst_r_sum2_0__0__q ;
wire Xd_0__inst_r_sum2_7__1__q ;
wire Xd_0__inst_r_sum2_6__1__q ;
wire Xd_0__inst_r_sum2_5__1__q ;
wire Xd_0__inst_r_sum2_4__1__q ;
wire Xd_0__inst_r_sum2_3__1__q ;
wire Xd_0__inst_r_sum2_2__1__q ;
wire Xd_0__inst_r_sum2_1__1__q ;
wire Xd_0__inst_r_sum2_0__1__q ;
wire Xd_0__inst_r_sum2_7__2__q ;
wire Xd_0__inst_r_sum2_6__2__q ;
wire Xd_0__inst_r_sum2_5__2__q ;
wire Xd_0__inst_r_sum2_4__2__q ;
wire Xd_0__inst_r_sum2_3__2__q ;
wire Xd_0__inst_r_sum2_2__2__q ;
wire Xd_0__inst_r_sum2_1__2__q ;
wire Xd_0__inst_r_sum2_0__2__q ;
wire Xd_0__inst_r_sum2_7__3__q ;
wire Xd_0__inst_r_sum2_6__3__q ;
wire Xd_0__inst_r_sum2_5__3__q ;
wire Xd_0__inst_r_sum2_4__3__q ;
wire Xd_0__inst_r_sum2_3__3__q ;
wire Xd_0__inst_r_sum2_2__3__q ;
wire Xd_0__inst_r_sum2_1__3__q ;
wire Xd_0__inst_r_sum2_0__3__q ;
wire Xd_0__inst_r_sum2_7__4__q ;
wire Xd_0__inst_r_sum2_6__4__q ;
wire Xd_0__inst_r_sum2_5__4__q ;
wire Xd_0__inst_r_sum2_4__4__q ;
wire Xd_0__inst_r_sum2_3__4__q ;
wire Xd_0__inst_r_sum2_2__4__q ;
wire Xd_0__inst_r_sum2_1__4__q ;
wire Xd_0__inst_r_sum2_0__4__q ;
wire Xd_0__inst_r_sum2_7__5__q ;
wire Xd_0__inst_r_sum2_6__5__q ;
wire Xd_0__inst_r_sum2_5__5__q ;
wire Xd_0__inst_r_sum2_4__5__q ;
wire Xd_0__inst_r_sum2_3__5__q ;
wire Xd_0__inst_r_sum2_2__5__q ;
wire Xd_0__inst_r_sum2_1__5__q ;
wire Xd_0__inst_r_sum2_0__5__q ;
wire Xd_0__inst_r_sum2_7__6__q ;
wire Xd_0__inst_r_sum2_6__6__q ;
wire Xd_0__inst_r_sum2_5__6__q ;
wire Xd_0__inst_r_sum2_4__6__q ;
wire Xd_0__inst_r_sum2_3__6__q ;
wire Xd_0__inst_r_sum2_2__6__q ;
wire Xd_0__inst_r_sum2_1__6__q ;
wire Xd_0__inst_r_sum2_0__6__q ;
wire Xd_0__inst_r_sum2_7__7__q ;
wire Xd_0__inst_r_sum2_6__7__q ;
wire Xd_0__inst_r_sum2_5__7__q ;
wire Xd_0__inst_r_sum2_4__7__q ;
wire Xd_0__inst_r_sum2_3__7__q ;
wire Xd_0__inst_r_sum2_2__7__q ;
wire Xd_0__inst_r_sum2_1__7__q ;
wire Xd_0__inst_r_sum2_0__7__q ;
wire Xd_0__inst_r_sum2_7__8__q ;
wire Xd_0__inst_r_sum2_6__8__q ;
wire Xd_0__inst_r_sum2_5__8__q ;
wire Xd_0__inst_r_sum2_4__8__q ;
wire Xd_0__inst_r_sum2_3__8__q ;
wire Xd_0__inst_r_sum2_2__8__q ;
wire Xd_0__inst_r_sum2_1__8__q ;
wire Xd_0__inst_r_sum2_0__8__q ;
wire Xd_0__inst_r_sum2_7__9__q ;
wire Xd_0__inst_r_sum2_6__9__q ;
wire Xd_0__inst_r_sum2_5__9__q ;
wire Xd_0__inst_r_sum2_4__9__q ;
wire Xd_0__inst_r_sum2_3__9__q ;
wire Xd_0__inst_r_sum2_2__9__q ;
wire Xd_0__inst_r_sum2_1__9__q ;
wire Xd_0__inst_r_sum2_0__9__q ;
wire Xd_0__inst_r_sum2_7__10__q ;
wire Xd_0__inst_r_sum2_6__10__q ;
wire Xd_0__inst_r_sum2_5__10__q ;
wire Xd_0__inst_r_sum2_4__10__q ;
wire Xd_0__inst_r_sum2_3__10__q ;
wire Xd_0__inst_r_sum2_2__10__q ;
wire Xd_0__inst_r_sum2_1__10__q ;
wire Xd_0__inst_r_sum2_0__10__q ;
wire Xd_0__inst_r_sum2_7__11__q ;
wire Xd_0__inst_r_sum2_6__11__q ;
wire Xd_0__inst_r_sum2_5__11__q ;
wire Xd_0__inst_r_sum2_4__11__q ;
wire Xd_0__inst_r_sum2_3__11__q ;
wire Xd_0__inst_r_sum2_2__11__q ;
wire Xd_0__inst_r_sum2_1__11__q ;
wire Xd_0__inst_r_sum2_0__11__q ;
wire Xd_0__inst_r_sum2_7__12__q ;
wire Xd_0__inst_r_sum2_6__12__q ;
wire Xd_0__inst_r_sum2_5__12__q ;
wire Xd_0__inst_r_sum2_4__12__q ;
wire Xd_0__inst_r_sum2_3__12__q ;
wire Xd_0__inst_r_sum2_2__12__q ;
wire Xd_0__inst_r_sum2_1__12__q ;
wire Xd_0__inst_r_sum2_0__12__q ;
wire Xd_0__inst_r_sum2_7__13__q ;
wire Xd_0__inst_r_sum2_6__13__q ;
wire Xd_0__inst_r_sum2_5__13__q ;
wire Xd_0__inst_r_sum2_4__13__q ;
wire Xd_0__inst_r_sum2_3__13__q ;
wire Xd_0__inst_r_sum2_2__13__q ;
wire Xd_0__inst_r_sum2_1__13__q ;
wire Xd_0__inst_r_sum2_0__13__q ;
wire Xd_0__inst_r_sum2_7__14__q ;
wire Xd_0__inst_r_sum2_6__14__q ;
wire Xd_0__inst_r_sum2_5__14__q ;
wire Xd_0__inst_r_sum2_4__14__q ;
wire Xd_0__inst_r_sum2_3__14__q ;
wire Xd_0__inst_r_sum2_2__14__q ;
wire Xd_0__inst_r_sum2_1__14__q ;
wire Xd_0__inst_r_sum2_0__14__q ;
wire Xd_0__inst_r_sum2_7__15__q ;
wire Xd_0__inst_r_sum2_6__15__q ;
wire Xd_0__inst_r_sum2_5__15__q ;
wire Xd_0__inst_r_sum2_4__15__q ;
wire Xd_0__inst_r_sum2_3__15__q ;
wire Xd_0__inst_r_sum2_2__15__q ;
wire Xd_0__inst_r_sum2_1__15__q ;
wire Xd_0__inst_r_sum2_0__15__q ;
wire Xd_0__inst_r_sum2_7__16__q ;
wire Xd_0__inst_r_sum2_6__16__q ;
wire Xd_0__inst_r_sum2_5__16__q ;
wire Xd_0__inst_r_sum2_4__16__q ;
wire Xd_0__inst_r_sum2_3__16__q ;
wire Xd_0__inst_r_sum2_2__16__q ;
wire Xd_0__inst_r_sum2_1__16__q ;
wire Xd_0__inst_r_sum2_0__16__q ;
wire Xd_0__inst_r_sum1_15__0__q ;
wire Xd_0__inst_r_sum1_14__0__q ;
wire Xd_0__inst_r_sum1_13__0__q ;
wire Xd_0__inst_r_sum1_12__0__q ;
wire Xd_0__inst_r_sum1_11__0__q ;
wire Xd_0__inst_r_sum1_10__0__q ;
wire Xd_0__inst_r_sum1_9__0__q ;
wire Xd_0__inst_r_sum1_8__0__q ;
wire Xd_0__inst_r_sum1_7__0__q ;
wire Xd_0__inst_r_sum1_6__0__q ;
wire Xd_0__inst_r_sum1_5__0__q ;
wire Xd_0__inst_r_sum1_4__0__q ;
wire Xd_0__inst_r_sum1_3__0__q ;
wire Xd_0__inst_r_sum1_2__0__q ;
wire Xd_0__inst_r_sum1_1__0__q ;
wire Xd_0__inst_r_sum1_0__0__q ;
wire Xd_0__inst_r_sum1_15__1__q ;
wire Xd_0__inst_r_sum1_14__1__q ;
wire Xd_0__inst_r_sum1_13__1__q ;
wire Xd_0__inst_r_sum1_12__1__q ;
wire Xd_0__inst_r_sum1_11__1__q ;
wire Xd_0__inst_r_sum1_10__1__q ;
wire Xd_0__inst_r_sum1_9__1__q ;
wire Xd_0__inst_r_sum1_8__1__q ;
wire Xd_0__inst_r_sum1_7__1__q ;
wire Xd_0__inst_r_sum1_6__1__q ;
wire Xd_0__inst_r_sum1_5__1__q ;
wire Xd_0__inst_r_sum1_4__1__q ;
wire Xd_0__inst_r_sum1_3__1__q ;
wire Xd_0__inst_r_sum1_2__1__q ;
wire Xd_0__inst_r_sum1_1__1__q ;
wire Xd_0__inst_r_sum1_0__1__q ;
wire Xd_0__inst_r_sum1_15__2__q ;
wire Xd_0__inst_r_sum1_14__2__q ;
wire Xd_0__inst_r_sum1_13__2__q ;
wire Xd_0__inst_r_sum1_12__2__q ;
wire Xd_0__inst_r_sum1_11__2__q ;
wire Xd_0__inst_r_sum1_10__2__q ;
wire Xd_0__inst_r_sum1_9__2__q ;
wire Xd_0__inst_r_sum1_8__2__q ;
wire Xd_0__inst_r_sum1_7__2__q ;
wire Xd_0__inst_r_sum1_6__2__q ;
wire Xd_0__inst_r_sum1_5__2__q ;
wire Xd_0__inst_r_sum1_4__2__q ;
wire Xd_0__inst_r_sum1_3__2__q ;
wire Xd_0__inst_r_sum1_2__2__q ;
wire Xd_0__inst_r_sum1_1__2__q ;
wire Xd_0__inst_r_sum1_0__2__q ;
wire Xd_0__inst_r_sum1_15__3__q ;
wire Xd_0__inst_r_sum1_14__3__q ;
wire Xd_0__inst_r_sum1_13__3__q ;
wire Xd_0__inst_r_sum1_12__3__q ;
wire Xd_0__inst_r_sum1_11__3__q ;
wire Xd_0__inst_r_sum1_10__3__q ;
wire Xd_0__inst_r_sum1_9__3__q ;
wire Xd_0__inst_r_sum1_8__3__q ;
wire Xd_0__inst_r_sum1_7__3__q ;
wire Xd_0__inst_r_sum1_6__3__q ;
wire Xd_0__inst_r_sum1_5__3__q ;
wire Xd_0__inst_r_sum1_4__3__q ;
wire Xd_0__inst_r_sum1_3__3__q ;
wire Xd_0__inst_r_sum1_2__3__q ;
wire Xd_0__inst_r_sum1_1__3__q ;
wire Xd_0__inst_r_sum1_0__3__q ;
wire Xd_0__inst_r_sum1_15__4__q ;
wire Xd_0__inst_r_sum1_14__4__q ;
wire Xd_0__inst_r_sum1_13__4__q ;
wire Xd_0__inst_r_sum1_12__4__q ;
wire Xd_0__inst_r_sum1_11__4__q ;
wire Xd_0__inst_r_sum1_10__4__q ;
wire Xd_0__inst_r_sum1_9__4__q ;
wire Xd_0__inst_r_sum1_8__4__q ;
wire Xd_0__inst_r_sum1_7__4__q ;
wire Xd_0__inst_r_sum1_6__4__q ;
wire Xd_0__inst_r_sum1_5__4__q ;
wire Xd_0__inst_r_sum1_4__4__q ;
wire Xd_0__inst_r_sum1_3__4__q ;
wire Xd_0__inst_r_sum1_2__4__q ;
wire Xd_0__inst_r_sum1_1__4__q ;
wire Xd_0__inst_r_sum1_0__4__q ;
wire Xd_0__inst_r_sum1_15__5__q ;
wire Xd_0__inst_r_sum1_14__5__q ;
wire Xd_0__inst_r_sum1_13__5__q ;
wire Xd_0__inst_r_sum1_12__5__q ;
wire Xd_0__inst_r_sum1_11__5__q ;
wire Xd_0__inst_r_sum1_10__5__q ;
wire Xd_0__inst_r_sum1_9__5__q ;
wire Xd_0__inst_r_sum1_8__5__q ;
wire Xd_0__inst_r_sum1_7__5__q ;
wire Xd_0__inst_r_sum1_6__5__q ;
wire Xd_0__inst_r_sum1_5__5__q ;
wire Xd_0__inst_r_sum1_4__5__q ;
wire Xd_0__inst_r_sum1_3__5__q ;
wire Xd_0__inst_r_sum1_2__5__q ;
wire Xd_0__inst_r_sum1_1__5__q ;
wire Xd_0__inst_r_sum1_0__5__q ;
wire Xd_0__inst_r_sum1_15__6__q ;
wire Xd_0__inst_r_sum1_14__6__q ;
wire Xd_0__inst_r_sum1_13__6__q ;
wire Xd_0__inst_r_sum1_12__6__q ;
wire Xd_0__inst_r_sum1_11__6__q ;
wire Xd_0__inst_r_sum1_10__6__q ;
wire Xd_0__inst_r_sum1_9__6__q ;
wire Xd_0__inst_r_sum1_8__6__q ;
wire Xd_0__inst_r_sum1_7__6__q ;
wire Xd_0__inst_r_sum1_6__6__q ;
wire Xd_0__inst_r_sum1_5__6__q ;
wire Xd_0__inst_r_sum1_4__6__q ;
wire Xd_0__inst_r_sum1_3__6__q ;
wire Xd_0__inst_r_sum1_2__6__q ;
wire Xd_0__inst_r_sum1_1__6__q ;
wire Xd_0__inst_r_sum1_0__6__q ;
wire Xd_0__inst_r_sum1_15__7__q ;
wire Xd_0__inst_r_sum1_14__7__q ;
wire Xd_0__inst_r_sum1_13__7__q ;
wire Xd_0__inst_r_sum1_12__7__q ;
wire Xd_0__inst_r_sum1_11__7__q ;
wire Xd_0__inst_r_sum1_10__7__q ;
wire Xd_0__inst_r_sum1_9__7__q ;
wire Xd_0__inst_r_sum1_8__7__q ;
wire Xd_0__inst_r_sum1_7__7__q ;
wire Xd_0__inst_r_sum1_6__7__q ;
wire Xd_0__inst_r_sum1_5__7__q ;
wire Xd_0__inst_r_sum1_4__7__q ;
wire Xd_0__inst_r_sum1_3__7__q ;
wire Xd_0__inst_r_sum1_2__7__q ;
wire Xd_0__inst_r_sum1_1__7__q ;
wire Xd_0__inst_r_sum1_0__7__q ;
wire Xd_0__inst_r_sum1_15__8__q ;
wire Xd_0__inst_r_sum1_14__8__q ;
wire Xd_0__inst_r_sum1_13__8__q ;
wire Xd_0__inst_r_sum1_12__8__q ;
wire Xd_0__inst_r_sum1_11__8__q ;
wire Xd_0__inst_r_sum1_10__8__q ;
wire Xd_0__inst_r_sum1_9__8__q ;
wire Xd_0__inst_r_sum1_8__8__q ;
wire Xd_0__inst_r_sum1_7__8__q ;
wire Xd_0__inst_r_sum1_6__8__q ;
wire Xd_0__inst_r_sum1_5__8__q ;
wire Xd_0__inst_r_sum1_4__8__q ;
wire Xd_0__inst_r_sum1_3__8__q ;
wire Xd_0__inst_r_sum1_2__8__q ;
wire Xd_0__inst_r_sum1_1__8__q ;
wire Xd_0__inst_r_sum1_0__8__q ;
wire Xd_0__inst_r_sum1_15__9__q ;
wire Xd_0__inst_r_sum1_14__9__q ;
wire Xd_0__inst_r_sum1_13__9__q ;
wire Xd_0__inst_r_sum1_12__9__q ;
wire Xd_0__inst_r_sum1_11__9__q ;
wire Xd_0__inst_r_sum1_10__9__q ;
wire Xd_0__inst_r_sum1_9__9__q ;
wire Xd_0__inst_r_sum1_8__9__q ;
wire Xd_0__inst_r_sum1_7__9__q ;
wire Xd_0__inst_r_sum1_6__9__q ;
wire Xd_0__inst_r_sum1_5__9__q ;
wire Xd_0__inst_r_sum1_4__9__q ;
wire Xd_0__inst_r_sum1_3__9__q ;
wire Xd_0__inst_r_sum1_2__9__q ;
wire Xd_0__inst_r_sum1_1__9__q ;
wire Xd_0__inst_r_sum1_0__9__q ;
wire Xd_0__inst_r_sum1_15__10__q ;
wire Xd_0__inst_r_sum1_14__10__q ;
wire Xd_0__inst_r_sum1_13__10__q ;
wire Xd_0__inst_r_sum1_12__10__q ;
wire Xd_0__inst_r_sum1_11__10__q ;
wire Xd_0__inst_r_sum1_10__10__q ;
wire Xd_0__inst_r_sum1_9__10__q ;
wire Xd_0__inst_r_sum1_8__10__q ;
wire Xd_0__inst_r_sum1_7__10__q ;
wire Xd_0__inst_r_sum1_6__10__q ;
wire Xd_0__inst_r_sum1_5__10__q ;
wire Xd_0__inst_r_sum1_4__10__q ;
wire Xd_0__inst_r_sum1_3__10__q ;
wire Xd_0__inst_r_sum1_2__10__q ;
wire Xd_0__inst_r_sum1_1__10__q ;
wire Xd_0__inst_r_sum1_0__10__q ;
wire Xd_0__inst_r_sum1_15__11__q ;
wire Xd_0__inst_r_sum1_14__11__q ;
wire Xd_0__inst_r_sum1_13__11__q ;
wire Xd_0__inst_r_sum1_12__11__q ;
wire Xd_0__inst_r_sum1_11__11__q ;
wire Xd_0__inst_r_sum1_10__11__q ;
wire Xd_0__inst_r_sum1_9__11__q ;
wire Xd_0__inst_r_sum1_8__11__q ;
wire Xd_0__inst_r_sum1_7__11__q ;
wire Xd_0__inst_r_sum1_6__11__q ;
wire Xd_0__inst_r_sum1_5__11__q ;
wire Xd_0__inst_r_sum1_4__11__q ;
wire Xd_0__inst_r_sum1_3__11__q ;
wire Xd_0__inst_r_sum1_2__11__q ;
wire Xd_0__inst_r_sum1_1__11__q ;
wire Xd_0__inst_r_sum1_0__11__q ;
wire Xd_0__inst_r_sum1_15__12__q ;
wire Xd_0__inst_r_sum1_14__12__q ;
wire Xd_0__inst_r_sum1_13__12__q ;
wire Xd_0__inst_r_sum1_12__12__q ;
wire Xd_0__inst_r_sum1_11__12__q ;
wire Xd_0__inst_r_sum1_10__12__q ;
wire Xd_0__inst_r_sum1_9__12__q ;
wire Xd_0__inst_r_sum1_8__12__q ;
wire Xd_0__inst_r_sum1_7__12__q ;
wire Xd_0__inst_r_sum1_6__12__q ;
wire Xd_0__inst_r_sum1_5__12__q ;
wire Xd_0__inst_r_sum1_4__12__q ;
wire Xd_0__inst_r_sum1_3__12__q ;
wire Xd_0__inst_r_sum1_2__12__q ;
wire Xd_0__inst_r_sum1_1__12__q ;
wire Xd_0__inst_r_sum1_0__12__q ;
wire Xd_0__inst_r_sum1_15__13__q ;
wire Xd_0__inst_r_sum1_14__13__q ;
wire Xd_0__inst_r_sum1_13__13__q ;
wire Xd_0__inst_r_sum1_12__13__q ;
wire Xd_0__inst_r_sum1_11__13__q ;
wire Xd_0__inst_r_sum1_10__13__q ;
wire Xd_0__inst_r_sum1_9__13__q ;
wire Xd_0__inst_r_sum1_8__13__q ;
wire Xd_0__inst_r_sum1_7__13__q ;
wire Xd_0__inst_r_sum1_6__13__q ;
wire Xd_0__inst_r_sum1_5__13__q ;
wire Xd_0__inst_r_sum1_4__13__q ;
wire Xd_0__inst_r_sum1_3__13__q ;
wire Xd_0__inst_r_sum1_2__13__q ;
wire Xd_0__inst_r_sum1_1__13__q ;
wire Xd_0__inst_r_sum1_0__13__q ;
wire Xd_0__inst_r_sum1_15__14__q ;
wire Xd_0__inst_r_sum1_14__14__q ;
wire Xd_0__inst_r_sum1_13__14__q ;
wire Xd_0__inst_r_sum1_12__14__q ;
wire Xd_0__inst_r_sum1_11__14__q ;
wire Xd_0__inst_r_sum1_10__14__q ;
wire Xd_0__inst_r_sum1_9__14__q ;
wire Xd_0__inst_r_sum1_8__14__q ;
wire Xd_0__inst_r_sum1_7__14__q ;
wire Xd_0__inst_r_sum1_6__14__q ;
wire Xd_0__inst_r_sum1_5__14__q ;
wire Xd_0__inst_r_sum1_4__14__q ;
wire Xd_0__inst_r_sum1_3__14__q ;
wire Xd_0__inst_r_sum1_2__14__q ;
wire Xd_0__inst_r_sum1_1__14__q ;
wire Xd_0__inst_r_sum1_0__14__q ;
wire Xd_0__inst_r_sum1_14__15__q ;
wire Xd_0__inst_r_sum1_15__15__q ;
wire Xd_0__inst_r_sum1_12__15__q ;
wire Xd_0__inst_r_sum1_13__15__q ;
wire Xd_0__inst_r_sum1_10__15__q ;
wire Xd_0__inst_r_sum1_11__15__q ;
wire Xd_0__inst_r_sum1_8__15__q ;
wire Xd_0__inst_r_sum1_9__15__q ;
wire Xd_0__inst_r_sum1_6__15__q ;
wire Xd_0__inst_r_sum1_7__15__q ;
wire Xd_0__inst_r_sum1_4__15__q ;
wire Xd_0__inst_r_sum1_5__15__q ;
wire Xd_0__inst_r_sum1_2__15__q ;
wire Xd_0__inst_r_sum1_3__15__q ;
wire Xd_0__inst_r_sum1_0__15__q ;
wire Xd_0__inst_r_sum1_1__15__q ;
wire Xd_0__inst_product_31__0__q ;
wire Xd_0__inst_product_30__0__q ;
wire Xd_0__inst_product_29__0__q ;
wire Xd_0__inst_product_28__0__q ;
wire Xd_0__inst_product_27__0__q ;
wire Xd_0__inst_product_26__0__q ;
wire Xd_0__inst_product_25__0__q ;
wire Xd_0__inst_product_24__0__q ;
wire Xd_0__inst_product_23__0__q ;
wire Xd_0__inst_product_22__0__q ;
wire Xd_0__inst_product_21__0__q ;
wire Xd_0__inst_product_20__0__q ;
wire Xd_0__inst_product_19__0__q ;
wire Xd_0__inst_product_18__0__q ;
wire Xd_0__inst_product_17__0__q ;
wire Xd_0__inst_product_16__0__q ;
wire Xd_0__inst_product_15__0__q ;
wire Xd_0__inst_product_14__0__q ;
wire Xd_0__inst_product_13__0__q ;
wire Xd_0__inst_product_12__0__q ;
wire Xd_0__inst_product_11__0__q ;
wire Xd_0__inst_product_10__0__q ;
wire Xd_0__inst_product_9__0__q ;
wire Xd_0__inst_product_8__0__q ;
wire Xd_0__inst_product_7__0__q ;
wire Xd_0__inst_product_6__0__q ;
wire Xd_0__inst_product_5__0__q ;
wire Xd_0__inst_product_4__0__q ;
wire Xd_0__inst_product_3__0__q ;
wire Xd_0__inst_product_2__0__q ;
wire Xd_0__inst_product_1__0__q ;
wire Xd_0__inst_product_0__0__q ;
wire Xd_0__inst_product_31__1__q ;
wire Xd_0__inst_product_30__1__q ;
wire Xd_0__inst_product_29__1__q ;
wire Xd_0__inst_product_28__1__q ;
wire Xd_0__inst_product_27__1__q ;
wire Xd_0__inst_product_26__1__q ;
wire Xd_0__inst_product_25__1__q ;
wire Xd_0__inst_product_24__1__q ;
wire Xd_0__inst_product_23__1__q ;
wire Xd_0__inst_product_22__1__q ;
wire Xd_0__inst_product_21__1__q ;
wire Xd_0__inst_product_20__1__q ;
wire Xd_0__inst_product_19__1__q ;
wire Xd_0__inst_product_18__1__q ;
wire Xd_0__inst_product_17__1__q ;
wire Xd_0__inst_product_16__1__q ;
wire Xd_0__inst_product_15__1__q ;
wire Xd_0__inst_product_14__1__q ;
wire Xd_0__inst_product_13__1__q ;
wire Xd_0__inst_product_12__1__q ;
wire Xd_0__inst_product_11__1__q ;
wire Xd_0__inst_product_10__1__q ;
wire Xd_0__inst_product_9__1__q ;
wire Xd_0__inst_product_8__1__q ;
wire Xd_0__inst_product_7__1__q ;
wire Xd_0__inst_product_6__1__q ;
wire Xd_0__inst_product_5__1__q ;
wire Xd_0__inst_product_4__1__q ;
wire Xd_0__inst_product_3__1__q ;
wire Xd_0__inst_product_2__1__q ;
wire Xd_0__inst_product_1__1__q ;
wire Xd_0__inst_product_0__1__q ;
wire Xd_0__inst_product_31__2__q ;
wire Xd_0__inst_product_30__2__q ;
wire Xd_0__inst_product_29__2__q ;
wire Xd_0__inst_product_28__2__q ;
wire Xd_0__inst_product_27__2__q ;
wire Xd_0__inst_product_26__2__q ;
wire Xd_0__inst_product_25__2__q ;
wire Xd_0__inst_product_24__2__q ;
wire Xd_0__inst_product_23__2__q ;
wire Xd_0__inst_product_22__2__q ;
wire Xd_0__inst_product_21__2__q ;
wire Xd_0__inst_product_20__2__q ;
wire Xd_0__inst_product_19__2__q ;
wire Xd_0__inst_product_18__2__q ;
wire Xd_0__inst_product_17__2__q ;
wire Xd_0__inst_product_16__2__q ;
wire Xd_0__inst_product_15__2__q ;
wire Xd_0__inst_product_14__2__q ;
wire Xd_0__inst_product_13__2__q ;
wire Xd_0__inst_product_12__2__q ;
wire Xd_0__inst_product_11__2__q ;
wire Xd_0__inst_product_10__2__q ;
wire Xd_0__inst_product_9__2__q ;
wire Xd_0__inst_product_8__2__q ;
wire Xd_0__inst_product_7__2__q ;
wire Xd_0__inst_product_6__2__q ;
wire Xd_0__inst_product_5__2__q ;
wire Xd_0__inst_product_4__2__q ;
wire Xd_0__inst_product_3__2__q ;
wire Xd_0__inst_product_2__2__q ;
wire Xd_0__inst_product_1__2__q ;
wire Xd_0__inst_product_0__2__q ;
wire Xd_0__inst_product_31__3__q ;
wire Xd_0__inst_product_30__3__q ;
wire Xd_0__inst_product_29__3__q ;
wire Xd_0__inst_product_28__3__q ;
wire Xd_0__inst_product_27__3__q ;
wire Xd_0__inst_product_26__3__q ;
wire Xd_0__inst_product_25__3__q ;
wire Xd_0__inst_product_24__3__q ;
wire Xd_0__inst_product_23__3__q ;
wire Xd_0__inst_product_22__3__q ;
wire Xd_0__inst_product_21__3__q ;
wire Xd_0__inst_product_20__3__q ;
wire Xd_0__inst_product_19__3__q ;
wire Xd_0__inst_product_18__3__q ;
wire Xd_0__inst_product_17__3__q ;
wire Xd_0__inst_product_16__3__q ;
wire Xd_0__inst_product_15__3__q ;
wire Xd_0__inst_product_14__3__q ;
wire Xd_0__inst_product_13__3__q ;
wire Xd_0__inst_product_12__3__q ;
wire Xd_0__inst_product_11__3__q ;
wire Xd_0__inst_product_10__3__q ;
wire Xd_0__inst_product_9__3__q ;
wire Xd_0__inst_product_8__3__q ;
wire Xd_0__inst_product_7__3__q ;
wire Xd_0__inst_product_6__3__q ;
wire Xd_0__inst_product_5__3__q ;
wire Xd_0__inst_product_4__3__q ;
wire Xd_0__inst_product_3__3__q ;
wire Xd_0__inst_product_2__3__q ;
wire Xd_0__inst_product_1__3__q ;
wire Xd_0__inst_product_0__3__q ;
wire Xd_0__inst_product_31__4__q ;
wire Xd_0__inst_product_30__4__q ;
wire Xd_0__inst_product_29__4__q ;
wire Xd_0__inst_product_28__4__q ;
wire Xd_0__inst_product_27__4__q ;
wire Xd_0__inst_product_26__4__q ;
wire Xd_0__inst_product_25__4__q ;
wire Xd_0__inst_product_24__4__q ;
wire Xd_0__inst_product_23__4__q ;
wire Xd_0__inst_product_22__4__q ;
wire Xd_0__inst_product_21__4__q ;
wire Xd_0__inst_product_20__4__q ;
wire Xd_0__inst_product_19__4__q ;
wire Xd_0__inst_product_18__4__q ;
wire Xd_0__inst_product_17__4__q ;
wire Xd_0__inst_product_16__4__q ;
wire Xd_0__inst_product_15__4__q ;
wire Xd_0__inst_product_14__4__q ;
wire Xd_0__inst_product_13__4__q ;
wire Xd_0__inst_product_12__4__q ;
wire Xd_0__inst_product_11__4__q ;
wire Xd_0__inst_product_10__4__q ;
wire Xd_0__inst_product_9__4__q ;
wire Xd_0__inst_product_8__4__q ;
wire Xd_0__inst_product_7__4__q ;
wire Xd_0__inst_product_6__4__q ;
wire Xd_0__inst_product_5__4__q ;
wire Xd_0__inst_product_4__4__q ;
wire Xd_0__inst_product_3__4__q ;
wire Xd_0__inst_product_2__4__q ;
wire Xd_0__inst_product_1__4__q ;
wire Xd_0__inst_product_0__4__q ;
wire Xd_0__inst_product_31__5__q ;
wire Xd_0__inst_product_30__5__q ;
wire Xd_0__inst_product_29__5__q ;
wire Xd_0__inst_product_28__5__q ;
wire Xd_0__inst_product_27__5__q ;
wire Xd_0__inst_product_26__5__q ;
wire Xd_0__inst_product_25__5__q ;
wire Xd_0__inst_product_24__5__q ;
wire Xd_0__inst_product_23__5__q ;
wire Xd_0__inst_product_22__5__q ;
wire Xd_0__inst_product_21__5__q ;
wire Xd_0__inst_product_20__5__q ;
wire Xd_0__inst_product_19__5__q ;
wire Xd_0__inst_product_18__5__q ;
wire Xd_0__inst_product_17__5__q ;
wire Xd_0__inst_product_16__5__q ;
wire Xd_0__inst_product_15__5__q ;
wire Xd_0__inst_product_14__5__q ;
wire Xd_0__inst_product_13__5__q ;
wire Xd_0__inst_product_12__5__q ;
wire Xd_0__inst_product_11__5__q ;
wire Xd_0__inst_product_10__5__q ;
wire Xd_0__inst_product_9__5__q ;
wire Xd_0__inst_product_8__5__q ;
wire Xd_0__inst_product_7__5__q ;
wire Xd_0__inst_product_6__5__q ;
wire Xd_0__inst_product_5__5__q ;
wire Xd_0__inst_product_4__5__q ;
wire Xd_0__inst_product_3__5__q ;
wire Xd_0__inst_product_2__5__q ;
wire Xd_0__inst_product_1__5__q ;
wire Xd_0__inst_product_0__5__q ;
wire Xd_0__inst_product_31__6__q ;
wire Xd_0__inst_product_30__6__q ;
wire Xd_0__inst_product_29__6__q ;
wire Xd_0__inst_product_28__6__q ;
wire Xd_0__inst_product_27__6__q ;
wire Xd_0__inst_product_26__6__q ;
wire Xd_0__inst_product_25__6__q ;
wire Xd_0__inst_product_24__6__q ;
wire Xd_0__inst_product_23__6__q ;
wire Xd_0__inst_product_22__6__q ;
wire Xd_0__inst_product_21__6__q ;
wire Xd_0__inst_product_20__6__q ;
wire Xd_0__inst_product_19__6__q ;
wire Xd_0__inst_product_18__6__q ;
wire Xd_0__inst_product_17__6__q ;
wire Xd_0__inst_product_16__6__q ;
wire Xd_0__inst_product_15__6__q ;
wire Xd_0__inst_product_14__6__q ;
wire Xd_0__inst_product_13__6__q ;
wire Xd_0__inst_product_12__6__q ;
wire Xd_0__inst_product_11__6__q ;
wire Xd_0__inst_product_10__6__q ;
wire Xd_0__inst_product_9__6__q ;
wire Xd_0__inst_product_8__6__q ;
wire Xd_0__inst_product_7__6__q ;
wire Xd_0__inst_product_6__6__q ;
wire Xd_0__inst_product_5__6__q ;
wire Xd_0__inst_product_4__6__q ;
wire Xd_0__inst_product_3__6__q ;
wire Xd_0__inst_product_2__6__q ;
wire Xd_0__inst_product_1__6__q ;
wire Xd_0__inst_product_0__6__q ;
wire Xd_0__inst_product_31__7__q ;
wire Xd_0__inst_product_30__7__q ;
wire Xd_0__inst_product_29__7__q ;
wire Xd_0__inst_product_28__7__q ;
wire Xd_0__inst_product_27__7__q ;
wire Xd_0__inst_product_26__7__q ;
wire Xd_0__inst_product_25__7__q ;
wire Xd_0__inst_product_24__7__q ;
wire Xd_0__inst_product_23__7__q ;
wire Xd_0__inst_product_22__7__q ;
wire Xd_0__inst_product_21__7__q ;
wire Xd_0__inst_product_20__7__q ;
wire Xd_0__inst_product_19__7__q ;
wire Xd_0__inst_product_18__7__q ;
wire Xd_0__inst_product_17__7__q ;
wire Xd_0__inst_product_16__7__q ;
wire Xd_0__inst_product_15__7__q ;
wire Xd_0__inst_product_14__7__q ;
wire Xd_0__inst_product_13__7__q ;
wire Xd_0__inst_product_12__7__q ;
wire Xd_0__inst_product_11__7__q ;
wire Xd_0__inst_product_10__7__q ;
wire Xd_0__inst_product_9__7__q ;
wire Xd_0__inst_product_8__7__q ;
wire Xd_0__inst_product_7__7__q ;
wire Xd_0__inst_product_6__7__q ;
wire Xd_0__inst_product_5__7__q ;
wire Xd_0__inst_product_4__7__q ;
wire Xd_0__inst_product_3__7__q ;
wire Xd_0__inst_product_2__7__q ;
wire Xd_0__inst_product_1__7__q ;
wire Xd_0__inst_product_0__7__q ;
wire Xd_0__inst_product_31__8__q ;
wire Xd_0__inst_product_30__8__q ;
wire Xd_0__inst_product_29__8__q ;
wire Xd_0__inst_product_28__8__q ;
wire Xd_0__inst_product_27__8__q ;
wire Xd_0__inst_product_26__8__q ;
wire Xd_0__inst_product_25__8__q ;
wire Xd_0__inst_product_24__8__q ;
wire Xd_0__inst_product_23__8__q ;
wire Xd_0__inst_product_22__8__q ;
wire Xd_0__inst_product_21__8__q ;
wire Xd_0__inst_product_20__8__q ;
wire Xd_0__inst_product_19__8__q ;
wire Xd_0__inst_product_18__8__q ;
wire Xd_0__inst_product_17__8__q ;
wire Xd_0__inst_product_16__8__q ;
wire Xd_0__inst_product_15__8__q ;
wire Xd_0__inst_product_14__8__q ;
wire Xd_0__inst_product_13__8__q ;
wire Xd_0__inst_product_12__8__q ;
wire Xd_0__inst_product_11__8__q ;
wire Xd_0__inst_product_10__8__q ;
wire Xd_0__inst_product_9__8__q ;
wire Xd_0__inst_product_8__8__q ;
wire Xd_0__inst_product_7__8__q ;
wire Xd_0__inst_product_6__8__q ;
wire Xd_0__inst_product_5__8__q ;
wire Xd_0__inst_product_4__8__q ;
wire Xd_0__inst_product_3__8__q ;
wire Xd_0__inst_product_2__8__q ;
wire Xd_0__inst_product_1__8__q ;
wire Xd_0__inst_product_0__8__q ;
wire Xd_0__inst_product_31__9__q ;
wire Xd_0__inst_product_30__9__q ;
wire Xd_0__inst_product_29__9__q ;
wire Xd_0__inst_product_28__9__q ;
wire Xd_0__inst_product_27__9__q ;
wire Xd_0__inst_product_26__9__q ;
wire Xd_0__inst_product_25__9__q ;
wire Xd_0__inst_product_24__9__q ;
wire Xd_0__inst_product_23__9__q ;
wire Xd_0__inst_product_22__9__q ;
wire Xd_0__inst_product_21__9__q ;
wire Xd_0__inst_product_20__9__q ;
wire Xd_0__inst_product_19__9__q ;
wire Xd_0__inst_product_18__9__q ;
wire Xd_0__inst_product_17__9__q ;
wire Xd_0__inst_product_16__9__q ;
wire Xd_0__inst_product_15__9__q ;
wire Xd_0__inst_product_14__9__q ;
wire Xd_0__inst_product_13__9__q ;
wire Xd_0__inst_product_12__9__q ;
wire Xd_0__inst_product_11__9__q ;
wire Xd_0__inst_product_10__9__q ;
wire Xd_0__inst_product_9__9__q ;
wire Xd_0__inst_product_8__9__q ;
wire Xd_0__inst_product_7__9__q ;
wire Xd_0__inst_product_6__9__q ;
wire Xd_0__inst_product_5__9__q ;
wire Xd_0__inst_product_4__9__q ;
wire Xd_0__inst_product_3__9__q ;
wire Xd_0__inst_product_2__9__q ;
wire Xd_0__inst_product_1__9__q ;
wire Xd_0__inst_product_0__9__q ;
wire Xd_0__inst_product_31__10__q ;
wire Xd_0__inst_product_30__10__q ;
wire Xd_0__inst_product_29__10__q ;
wire Xd_0__inst_product_28__10__q ;
wire Xd_0__inst_product_27__10__q ;
wire Xd_0__inst_product_26__10__q ;
wire Xd_0__inst_product_25__10__q ;
wire Xd_0__inst_product_24__10__q ;
wire Xd_0__inst_product_23__10__q ;
wire Xd_0__inst_product_22__10__q ;
wire Xd_0__inst_product_21__10__q ;
wire Xd_0__inst_product_20__10__q ;
wire Xd_0__inst_product_19__10__q ;
wire Xd_0__inst_product_18__10__q ;
wire Xd_0__inst_product_17__10__q ;
wire Xd_0__inst_product_16__10__q ;
wire Xd_0__inst_product_15__10__q ;
wire Xd_0__inst_product_14__10__q ;
wire Xd_0__inst_product_13__10__q ;
wire Xd_0__inst_product_12__10__q ;
wire Xd_0__inst_product_11__10__q ;
wire Xd_0__inst_product_10__10__q ;
wire Xd_0__inst_product_9__10__q ;
wire Xd_0__inst_product_8__10__q ;
wire Xd_0__inst_product_7__10__q ;
wire Xd_0__inst_product_6__10__q ;
wire Xd_0__inst_product_5__10__q ;
wire Xd_0__inst_product_4__10__q ;
wire Xd_0__inst_product_3__10__q ;
wire Xd_0__inst_product_2__10__q ;
wire Xd_0__inst_product_1__10__q ;
wire Xd_0__inst_product_0__10__q ;
wire Xd_0__inst_product_31__11__q ;
wire Xd_0__inst_product_30__11__q ;
wire Xd_0__inst_product_29__11__q ;
wire Xd_0__inst_product_28__11__q ;
wire Xd_0__inst_product_27__11__q ;
wire Xd_0__inst_product_26__11__q ;
wire Xd_0__inst_product_25__11__q ;
wire Xd_0__inst_product_24__11__q ;
wire Xd_0__inst_product_23__11__q ;
wire Xd_0__inst_product_22__11__q ;
wire Xd_0__inst_product_21__11__q ;
wire Xd_0__inst_product_20__11__q ;
wire Xd_0__inst_product_19__11__q ;
wire Xd_0__inst_product_18__11__q ;
wire Xd_0__inst_product_17__11__q ;
wire Xd_0__inst_product_16__11__q ;
wire Xd_0__inst_product_15__11__q ;
wire Xd_0__inst_product_14__11__q ;
wire Xd_0__inst_product_13__11__q ;
wire Xd_0__inst_product_12__11__q ;
wire Xd_0__inst_product_11__11__q ;
wire Xd_0__inst_product_10__11__q ;
wire Xd_0__inst_product_9__11__q ;
wire Xd_0__inst_product_8__11__q ;
wire Xd_0__inst_product_7__11__q ;
wire Xd_0__inst_product_6__11__q ;
wire Xd_0__inst_product_5__11__q ;
wire Xd_0__inst_product_4__11__q ;
wire Xd_0__inst_product_3__11__q ;
wire Xd_0__inst_product_2__11__q ;
wire Xd_0__inst_product_1__11__q ;
wire Xd_0__inst_product_0__11__q ;
wire Xd_0__inst_product_31__12__q ;
wire Xd_0__inst_product_30__12__q ;
wire Xd_0__inst_product_29__12__q ;
wire Xd_0__inst_product_28__12__q ;
wire Xd_0__inst_product_27__12__q ;
wire Xd_0__inst_product_26__12__q ;
wire Xd_0__inst_product_25__12__q ;
wire Xd_0__inst_product_24__12__q ;
wire Xd_0__inst_product_23__12__q ;
wire Xd_0__inst_product_22__12__q ;
wire Xd_0__inst_product_21__12__q ;
wire Xd_0__inst_product_20__12__q ;
wire Xd_0__inst_product_19__12__q ;
wire Xd_0__inst_product_18__12__q ;
wire Xd_0__inst_product_17__12__q ;
wire Xd_0__inst_product_16__12__q ;
wire Xd_0__inst_product_15__12__q ;
wire Xd_0__inst_product_14__12__q ;
wire Xd_0__inst_product_13__12__q ;
wire Xd_0__inst_product_12__12__q ;
wire Xd_0__inst_product_11__12__q ;
wire Xd_0__inst_product_10__12__q ;
wire Xd_0__inst_product_9__12__q ;
wire Xd_0__inst_product_8__12__q ;
wire Xd_0__inst_product_7__12__q ;
wire Xd_0__inst_product_6__12__q ;
wire Xd_0__inst_product_5__12__q ;
wire Xd_0__inst_product_4__12__q ;
wire Xd_0__inst_product_3__12__q ;
wire Xd_0__inst_product_2__12__q ;
wire Xd_0__inst_product_1__12__q ;
wire Xd_0__inst_product_0__12__q ;
wire Xd_0__inst_product_31__13__q ;
wire Xd_0__inst_product_30__13__q ;
wire Xd_0__inst_product_29__13__q ;
wire Xd_0__inst_product_28__13__q ;
wire Xd_0__inst_product_27__13__q ;
wire Xd_0__inst_product_26__13__q ;
wire Xd_0__inst_product_25__13__q ;
wire Xd_0__inst_product_24__13__q ;
wire Xd_0__inst_product_23__13__q ;
wire Xd_0__inst_product_22__13__q ;
wire Xd_0__inst_product_21__13__q ;
wire Xd_0__inst_product_20__13__q ;
wire Xd_0__inst_product_19__13__q ;
wire Xd_0__inst_product_18__13__q ;
wire Xd_0__inst_product_17__13__q ;
wire Xd_0__inst_product_16__13__q ;
wire Xd_0__inst_product_15__13__q ;
wire Xd_0__inst_product_14__13__q ;
wire Xd_0__inst_product_13__13__q ;
wire Xd_0__inst_product_12__13__q ;
wire Xd_0__inst_product_11__13__q ;
wire Xd_0__inst_product_10__13__q ;
wire Xd_0__inst_product_9__13__q ;
wire Xd_0__inst_product_8__13__q ;
wire Xd_0__inst_product_7__13__q ;
wire Xd_0__inst_product_6__13__q ;
wire Xd_0__inst_product_5__13__q ;
wire Xd_0__inst_product_4__13__q ;
wire Xd_0__inst_product_3__13__q ;
wire Xd_0__inst_product_2__13__q ;
wire Xd_0__inst_product_1__13__q ;
wire Xd_0__inst_product_0__13__q ;
wire Xd_0__inst_product1_31__0__q ;
wire Xd_0__inst_product1_30__0__q ;
wire Xd_0__inst_product1_29__0__q ;
wire Xd_0__inst_product1_28__0__q ;
wire Xd_0__inst_product1_27__0__q ;
wire Xd_0__inst_product1_26__0__q ;
wire Xd_0__inst_product1_25__0__q ;
wire Xd_0__inst_product1_24__0__q ;
wire Xd_0__inst_product1_23__0__q ;
wire Xd_0__inst_product1_22__0__q ;
wire Xd_0__inst_product1_21__0__q ;
wire Xd_0__inst_product1_20__0__q ;
wire Xd_0__inst_product1_19__0__q ;
wire Xd_0__inst_product1_18__0__q ;
wire Xd_0__inst_product1_17__0__q ;
wire Xd_0__inst_product1_16__0__q ;
wire Xd_0__inst_product1_15__0__q ;
wire Xd_0__inst_product1_14__0__q ;
wire Xd_0__inst_product1_13__0__q ;
wire Xd_0__inst_product1_12__0__q ;
wire Xd_0__inst_product1_11__0__q ;
wire Xd_0__inst_product1_10__0__q ;
wire Xd_0__inst_product1_9__0__q ;
wire Xd_0__inst_product1_8__0__q ;
wire Xd_0__inst_product1_7__0__q ;
wire Xd_0__inst_product1_6__0__q ;
wire Xd_0__inst_product1_5__0__q ;
wire Xd_0__inst_product1_4__0__q ;
wire Xd_0__inst_product1_3__0__q ;
wire Xd_0__inst_product1_2__0__q ;
wire Xd_0__inst_product1_1__0__q ;
wire Xd_0__inst_product1_0__0__q ;
wire Xd_0__inst_product1_31__1__q ;
wire Xd_0__inst_product1_30__1__q ;
wire Xd_0__inst_product1_29__1__q ;
wire Xd_0__inst_product1_28__1__q ;
wire Xd_0__inst_product1_27__1__q ;
wire Xd_0__inst_product1_26__1__q ;
wire Xd_0__inst_product1_25__1__q ;
wire Xd_0__inst_product1_24__1__q ;
wire Xd_0__inst_product1_23__1__q ;
wire Xd_0__inst_product1_22__1__q ;
wire Xd_0__inst_product1_21__1__q ;
wire Xd_0__inst_product1_20__1__q ;
wire Xd_0__inst_product1_19__1__q ;
wire Xd_0__inst_product1_18__1__q ;
wire Xd_0__inst_product1_17__1__q ;
wire Xd_0__inst_product1_16__1__q ;
wire Xd_0__inst_product1_15__1__q ;
wire Xd_0__inst_product1_14__1__q ;
wire Xd_0__inst_product1_13__1__q ;
wire Xd_0__inst_product1_12__1__q ;
wire Xd_0__inst_product1_11__1__q ;
wire Xd_0__inst_product1_10__1__q ;
wire Xd_0__inst_product1_9__1__q ;
wire Xd_0__inst_product1_8__1__q ;
wire Xd_0__inst_product1_7__1__q ;
wire Xd_0__inst_product1_6__1__q ;
wire Xd_0__inst_product1_5__1__q ;
wire Xd_0__inst_product1_4__1__q ;
wire Xd_0__inst_product1_3__1__q ;
wire Xd_0__inst_product1_2__1__q ;
wire Xd_0__inst_product1_1__1__q ;
wire Xd_0__inst_product1_0__1__q ;
wire Xd_0__inst_product1_31__2__q ;
wire Xd_0__inst_product1_30__2__q ;
wire Xd_0__inst_product1_29__2__q ;
wire Xd_0__inst_product1_28__2__q ;
wire Xd_0__inst_product1_27__2__q ;
wire Xd_0__inst_product1_26__2__q ;
wire Xd_0__inst_product1_25__2__q ;
wire Xd_0__inst_product1_24__2__q ;
wire Xd_0__inst_product1_23__2__q ;
wire Xd_0__inst_product1_22__2__q ;
wire Xd_0__inst_product1_21__2__q ;
wire Xd_0__inst_product1_20__2__q ;
wire Xd_0__inst_product1_19__2__q ;
wire Xd_0__inst_product1_18__2__q ;
wire Xd_0__inst_product1_17__2__q ;
wire Xd_0__inst_product1_16__2__q ;
wire Xd_0__inst_product1_15__2__q ;
wire Xd_0__inst_product1_14__2__q ;
wire Xd_0__inst_product1_13__2__q ;
wire Xd_0__inst_product1_12__2__q ;
wire Xd_0__inst_product1_11__2__q ;
wire Xd_0__inst_product1_10__2__q ;
wire Xd_0__inst_product1_9__2__q ;
wire Xd_0__inst_product1_8__2__q ;
wire Xd_0__inst_product1_7__2__q ;
wire Xd_0__inst_product1_6__2__q ;
wire Xd_0__inst_product1_5__2__q ;
wire Xd_0__inst_product1_4__2__q ;
wire Xd_0__inst_product1_3__2__q ;
wire Xd_0__inst_product1_2__2__q ;
wire Xd_0__inst_product1_1__2__q ;
wire Xd_0__inst_product1_0__2__q ;
wire Xd_0__inst_mult_31_0_q ;
wire Xd_0__inst_mult_31_1_q ;
wire Xd_0__inst_mult_30_0_q ;
wire Xd_0__inst_mult_30_1_q ;
wire Xd_0__inst_mult_29_0_q ;
wire Xd_0__inst_mult_29_1_q ;
wire Xd_0__inst_mult_28_0_q ;
wire Xd_0__inst_mult_28_1_q ;
wire Xd_0__inst_mult_27_0_q ;
wire Xd_0__inst_mult_27_1_q ;
wire Xd_0__inst_mult_26_0_q ;
wire Xd_0__inst_mult_26_1_q ;
wire Xd_0__inst_mult_25_0_q ;
wire Xd_0__inst_mult_25_1_q ;
wire Xd_0__inst_mult_24_0_q ;
wire Xd_0__inst_mult_24_1_q ;
wire Xd_0__inst_mult_23_0_q ;
wire Xd_0__inst_mult_23_1_q ;
wire Xd_0__inst_mult_22_0_q ;
wire Xd_0__inst_mult_22_1_q ;
wire Xd_0__inst_mult_21_0_q ;
wire Xd_0__inst_mult_21_1_q ;
wire Xd_0__inst_mult_20_0_q ;
wire Xd_0__inst_mult_20_1_q ;
wire Xd_0__inst_mult_19_0_q ;
wire Xd_0__inst_mult_19_1_q ;
wire Xd_0__inst_mult_18_0_q ;
wire Xd_0__inst_mult_18_1_q ;
wire Xd_0__inst_mult_17_0_q ;
wire Xd_0__inst_mult_17_1_q ;
wire Xd_0__inst_mult_16_0_q ;
wire Xd_0__inst_mult_16_1_q ;
wire Xd_0__inst_mult_15_0_q ;
wire Xd_0__inst_mult_15_1_q ;
wire Xd_0__inst_mult_14_0_q ;
wire Xd_0__inst_mult_14_1_q ;
wire Xd_0__inst_mult_13_0_q ;
wire Xd_0__inst_mult_13_1_q ;
wire Xd_0__inst_mult_12_0_q ;
wire Xd_0__inst_mult_12_1_q ;
wire Xd_0__inst_mult_11_0_q ;
wire Xd_0__inst_mult_11_1_q ;
wire Xd_0__inst_mult_10_0_q ;
wire Xd_0__inst_mult_10_1_q ;
wire Xd_0__inst_mult_9_0_q ;
wire Xd_0__inst_mult_9_1_q ;
wire Xd_0__inst_mult_8_0_q ;
wire Xd_0__inst_mult_8_1_q ;
wire Xd_0__inst_mult_7_0_q ;
wire Xd_0__inst_mult_7_1_q ;
wire Xd_0__inst_mult_6_0_q ;
wire Xd_0__inst_mult_6_1_q ;
wire Xd_0__inst_mult_5_0_q ;
wire Xd_0__inst_mult_5_1_q ;
wire Xd_0__inst_mult_4_0_q ;
wire Xd_0__inst_mult_4_1_q ;
wire Xd_0__inst_mult_3_0_q ;
wire Xd_0__inst_mult_3_1_q ;
wire Xd_0__inst_mult_2_0_q ;
wire Xd_0__inst_mult_2_1_q ;
wire Xd_0__inst_mult_1_0_q ;
wire Xd_0__inst_mult_1_1_q ;
wire Xd_0__inst_mult_0_0_q ;
wire Xd_0__inst_mult_0_1_q ;
wire Xd_0__inst_mult_31_2_q ;
wire Xd_0__inst_mult_31_3_q ;
wire Xd_0__inst_mult_30_2_q ;
wire Xd_0__inst_mult_30_3_q ;
wire Xd_0__inst_mult_29_2_q ;
wire Xd_0__inst_mult_29_3_q ;
wire Xd_0__inst_mult_28_2_q ;
wire Xd_0__inst_mult_28_3_q ;
wire Xd_0__inst_mult_27_2_q ;
wire Xd_0__inst_mult_27_3_q ;
wire Xd_0__inst_mult_26_2_q ;
wire Xd_0__inst_mult_26_3_q ;
wire Xd_0__inst_mult_25_2_q ;
wire Xd_0__inst_mult_25_3_q ;
wire Xd_0__inst_mult_24_2_q ;
wire Xd_0__inst_mult_24_3_q ;
wire Xd_0__inst_mult_23_2_q ;
wire Xd_0__inst_mult_23_3_q ;
wire Xd_0__inst_mult_22_2_q ;
wire Xd_0__inst_mult_22_3_q ;
wire Xd_0__inst_mult_21_2_q ;
wire Xd_0__inst_mult_21_3_q ;
wire Xd_0__inst_mult_20_2_q ;
wire Xd_0__inst_mult_20_3_q ;
wire Xd_0__inst_mult_19_2_q ;
wire Xd_0__inst_mult_19_3_q ;
wire Xd_0__inst_mult_18_2_q ;
wire Xd_0__inst_mult_18_3_q ;
wire Xd_0__inst_mult_17_2_q ;
wire Xd_0__inst_mult_17_3_q ;
wire Xd_0__inst_mult_16_2_q ;
wire Xd_0__inst_mult_16_3_q ;
wire Xd_0__inst_mult_15_2_q ;
wire Xd_0__inst_mult_15_3_q ;
wire Xd_0__inst_mult_14_2_q ;
wire Xd_0__inst_mult_14_3_q ;
wire Xd_0__inst_mult_13_2_q ;
wire Xd_0__inst_mult_13_3_q ;
wire Xd_0__inst_mult_12_2_q ;
wire Xd_0__inst_mult_12_3_q ;
wire Xd_0__inst_mult_11_2_q ;
wire Xd_0__inst_mult_11_3_q ;
wire Xd_0__inst_mult_10_2_q ;
wire Xd_0__inst_mult_10_3_q ;
wire Xd_0__inst_mult_9_2_q ;
wire Xd_0__inst_mult_9_3_q ;
wire Xd_0__inst_mult_8_2_q ;
wire Xd_0__inst_mult_8_3_q ;
wire Xd_0__inst_mult_7_2_q ;
wire Xd_0__inst_mult_7_3_q ;
wire Xd_0__inst_mult_6_2_q ;
wire Xd_0__inst_mult_6_3_q ;
wire Xd_0__inst_mult_5_2_q ;
wire Xd_0__inst_mult_5_3_q ;
wire Xd_0__inst_mult_4_2_q ;
wire Xd_0__inst_mult_4_3_q ;
wire Xd_0__inst_mult_3_2_q ;
wire Xd_0__inst_mult_3_3_q ;
wire Xd_0__inst_mult_2_2_q ;
wire Xd_0__inst_mult_2_3_q ;
wire Xd_0__inst_mult_1_2_q ;
wire Xd_0__inst_mult_1_3_q ;
wire Xd_0__inst_mult_0_2_q ;
wire Xd_0__inst_mult_0_3_q ;
wire Xd_0__inst_mult_31_4_q ;
wire Xd_0__inst_mult_31_5_q ;
wire Xd_0__inst_mult_30_4_q ;
wire Xd_0__inst_mult_30_5_q ;
wire Xd_0__inst_mult_29_4_q ;
wire Xd_0__inst_mult_29_5_q ;
wire Xd_0__inst_mult_28_4_q ;
wire Xd_0__inst_mult_28_5_q ;
wire Xd_0__inst_mult_27_4_q ;
wire Xd_0__inst_mult_27_5_q ;
wire Xd_0__inst_mult_26_4_q ;
wire Xd_0__inst_mult_26_5_q ;
wire Xd_0__inst_mult_25_4_q ;
wire Xd_0__inst_mult_25_5_q ;
wire Xd_0__inst_mult_24_4_q ;
wire Xd_0__inst_mult_24_5_q ;
wire Xd_0__inst_mult_23_4_q ;
wire Xd_0__inst_mult_23_5_q ;
wire Xd_0__inst_mult_22_4_q ;
wire Xd_0__inst_mult_22_5_q ;
wire Xd_0__inst_mult_21_4_q ;
wire Xd_0__inst_mult_21_5_q ;
wire Xd_0__inst_mult_20_4_q ;
wire Xd_0__inst_mult_20_5_q ;
wire Xd_0__inst_mult_19_4_q ;
wire Xd_0__inst_mult_19_5_q ;
wire Xd_0__inst_mult_18_4_q ;
wire Xd_0__inst_mult_18_5_q ;
wire Xd_0__inst_mult_17_4_q ;
wire Xd_0__inst_mult_17_5_q ;
wire Xd_0__inst_mult_16_4_q ;
wire Xd_0__inst_mult_16_5_q ;
wire Xd_0__inst_mult_15_4_q ;
wire Xd_0__inst_mult_15_5_q ;
wire Xd_0__inst_mult_14_4_q ;
wire Xd_0__inst_mult_14_5_q ;
wire Xd_0__inst_mult_13_4_q ;
wire Xd_0__inst_mult_13_5_q ;
wire Xd_0__inst_mult_12_4_q ;
wire Xd_0__inst_mult_12_5_q ;
wire Xd_0__inst_mult_11_4_q ;
wire Xd_0__inst_mult_11_5_q ;
wire Xd_0__inst_mult_10_4_q ;
wire Xd_0__inst_mult_10_5_q ;
wire Xd_0__inst_mult_9_4_q ;
wire Xd_0__inst_mult_9_5_q ;
wire Xd_0__inst_mult_8_4_q ;
wire Xd_0__inst_mult_8_5_q ;
wire Xd_0__inst_mult_7_4_q ;
wire Xd_0__inst_mult_7_5_q ;
wire Xd_0__inst_mult_6_4_q ;
wire Xd_0__inst_mult_6_5_q ;
wire Xd_0__inst_mult_5_4_q ;
wire Xd_0__inst_mult_5_5_q ;
wire Xd_0__inst_mult_4_4_q ;
wire Xd_0__inst_mult_4_5_q ;
wire Xd_0__inst_mult_3_4_q ;
wire Xd_0__inst_mult_3_5_q ;
wire Xd_0__inst_mult_2_4_q ;
wire Xd_0__inst_mult_2_5_q ;
wire Xd_0__inst_mult_1_4_q ;
wire Xd_0__inst_mult_1_5_q ;
wire Xd_0__inst_mult_0_4_q ;
wire Xd_0__inst_mult_0_5_q ;
wire Xd_0__inst_mult_31_6_q ;
wire Xd_0__inst_mult_31_7_q ;
wire Xd_0__inst_mult_30_6_q ;
wire Xd_0__inst_mult_30_7_q ;
wire Xd_0__inst_mult_29_6_q ;
wire Xd_0__inst_mult_29_7_q ;
wire Xd_0__inst_mult_28_6_q ;
wire Xd_0__inst_mult_28_7_q ;
wire Xd_0__inst_mult_27_6_q ;
wire Xd_0__inst_mult_27_7_q ;
wire Xd_0__inst_mult_26_6_q ;
wire Xd_0__inst_mult_26_7_q ;
wire Xd_0__inst_mult_25_6_q ;
wire Xd_0__inst_mult_25_7_q ;
wire Xd_0__inst_mult_24_6_q ;
wire Xd_0__inst_mult_24_7_q ;
wire Xd_0__inst_mult_23_6_q ;
wire Xd_0__inst_mult_23_7_q ;
wire Xd_0__inst_mult_22_6_q ;
wire Xd_0__inst_mult_22_7_q ;
wire Xd_0__inst_mult_21_6_q ;
wire Xd_0__inst_mult_21_7_q ;
wire Xd_0__inst_mult_20_6_q ;
wire Xd_0__inst_mult_20_7_q ;
wire Xd_0__inst_mult_19_6_q ;
wire Xd_0__inst_mult_19_7_q ;
wire Xd_0__inst_mult_18_6_q ;
wire Xd_0__inst_mult_18_7_q ;
wire Xd_0__inst_mult_17_6_q ;
wire Xd_0__inst_mult_17_7_q ;
wire Xd_0__inst_mult_16_6_q ;
wire Xd_0__inst_mult_16_7_q ;
wire Xd_0__inst_mult_15_6_q ;
wire Xd_0__inst_mult_15_7_q ;
wire Xd_0__inst_mult_14_6_q ;
wire Xd_0__inst_mult_14_7_q ;
wire Xd_0__inst_mult_13_6_q ;
wire Xd_0__inst_mult_13_7_q ;
wire Xd_0__inst_mult_12_6_q ;
wire Xd_0__inst_mult_12_7_q ;
wire Xd_0__inst_mult_11_6_q ;
wire Xd_0__inst_mult_11_7_q ;
wire Xd_0__inst_mult_10_6_q ;
wire Xd_0__inst_mult_10_7_q ;
wire Xd_0__inst_mult_9_6_q ;
wire Xd_0__inst_mult_9_7_q ;
wire Xd_0__inst_mult_8_6_q ;
wire Xd_0__inst_mult_8_7_q ;
wire Xd_0__inst_mult_7_6_q ;
wire Xd_0__inst_mult_7_7_q ;
wire Xd_0__inst_mult_6_6_q ;
wire Xd_0__inst_mult_6_7_q ;
wire Xd_0__inst_mult_5_6_q ;
wire Xd_0__inst_mult_5_7_q ;
wire Xd_0__inst_mult_4_6_q ;
wire Xd_0__inst_mult_4_7_q ;
wire Xd_0__inst_mult_3_6_q ;
wire Xd_0__inst_mult_3_7_q ;
wire Xd_0__inst_mult_2_6_q ;
wire Xd_0__inst_mult_2_7_q ;
wire Xd_0__inst_mult_1_6_q ;
wire Xd_0__inst_mult_1_7_q ;
wire Xd_0__inst_mult_0_6_q ;
wire Xd_0__inst_mult_0_7_q ;
wire Xd_0__inst_mult_31_8_q ;
wire Xd_0__inst_mult_31_9_q ;
wire Xd_0__inst_mult_30_8_q ;
wire Xd_0__inst_mult_30_9_q ;
wire Xd_0__inst_mult_29_8_q ;
wire Xd_0__inst_mult_29_9_q ;
wire Xd_0__inst_mult_28_8_q ;
wire Xd_0__inst_mult_28_9_q ;
wire Xd_0__inst_mult_27_8_q ;
wire Xd_0__inst_mult_27_9_q ;
wire Xd_0__inst_mult_26_8_q ;
wire Xd_0__inst_mult_26_9_q ;
wire Xd_0__inst_mult_25_8_q ;
wire Xd_0__inst_mult_25_9_q ;
wire Xd_0__inst_mult_24_8_q ;
wire Xd_0__inst_mult_24_9_q ;
wire Xd_0__inst_mult_23_8_q ;
wire Xd_0__inst_mult_23_9_q ;
wire Xd_0__inst_mult_22_8_q ;
wire Xd_0__inst_mult_22_9_q ;
wire Xd_0__inst_mult_21_8_q ;
wire Xd_0__inst_mult_21_9_q ;
wire Xd_0__inst_mult_20_8_q ;
wire Xd_0__inst_mult_20_9_q ;
wire Xd_0__inst_mult_19_8_q ;
wire Xd_0__inst_mult_19_9_q ;
wire Xd_0__inst_mult_18_8_q ;
wire Xd_0__inst_mult_18_9_q ;
wire Xd_0__inst_mult_17_8_q ;
wire Xd_0__inst_mult_17_9_q ;
wire Xd_0__inst_mult_16_8_q ;
wire Xd_0__inst_mult_16_9_q ;
wire Xd_0__inst_mult_15_8_q ;
wire Xd_0__inst_mult_15_9_q ;
wire Xd_0__inst_mult_14_8_q ;
wire Xd_0__inst_mult_14_9_q ;
wire Xd_0__inst_mult_13_8_q ;
wire Xd_0__inst_mult_13_9_q ;
wire Xd_0__inst_mult_12_8_q ;
wire Xd_0__inst_mult_12_9_q ;
wire Xd_0__inst_mult_11_8_q ;
wire Xd_0__inst_mult_11_9_q ;
wire Xd_0__inst_mult_10_8_q ;
wire Xd_0__inst_mult_10_9_q ;
wire Xd_0__inst_mult_9_8_q ;
wire Xd_0__inst_mult_9_9_q ;
wire Xd_0__inst_mult_8_8_q ;
wire Xd_0__inst_mult_8_9_q ;
wire Xd_0__inst_mult_7_8_q ;
wire Xd_0__inst_mult_7_9_q ;
wire Xd_0__inst_mult_6_8_q ;
wire Xd_0__inst_mult_6_9_q ;
wire Xd_0__inst_mult_5_8_q ;
wire Xd_0__inst_mult_5_9_q ;
wire Xd_0__inst_mult_4_8_q ;
wire Xd_0__inst_mult_4_9_q ;
wire Xd_0__inst_mult_3_8_q ;
wire Xd_0__inst_mult_3_9_q ;
wire Xd_0__inst_mult_2_8_q ;
wire Xd_0__inst_mult_2_9_q ;
wire Xd_0__inst_mult_1_8_q ;
wire Xd_0__inst_mult_1_9_q ;
wire Xd_0__inst_mult_0_8_q ;
wire Xd_0__inst_mult_0_9_q ;
wire Xd_0__inst_mult_31_10_q ;
wire Xd_0__inst_mult_31_11_q ;
wire Xd_0__inst_mult_30_10_q ;
wire Xd_0__inst_mult_30_11_q ;
wire Xd_0__inst_mult_29_10_q ;
wire Xd_0__inst_mult_29_11_q ;
wire Xd_0__inst_mult_28_10_q ;
wire Xd_0__inst_mult_28_11_q ;
wire Xd_0__inst_mult_27_10_q ;
wire Xd_0__inst_mult_27_11_q ;
wire Xd_0__inst_mult_26_10_q ;
wire Xd_0__inst_mult_26_11_q ;
wire Xd_0__inst_mult_25_10_q ;
wire Xd_0__inst_mult_25_11_q ;
wire Xd_0__inst_mult_24_10_q ;
wire Xd_0__inst_mult_24_11_q ;
wire Xd_0__inst_mult_23_10_q ;
wire Xd_0__inst_mult_23_11_q ;
wire Xd_0__inst_mult_22_10_q ;
wire Xd_0__inst_mult_22_11_q ;
wire Xd_0__inst_mult_21_10_q ;
wire Xd_0__inst_mult_21_11_q ;
wire Xd_0__inst_mult_20_10_q ;
wire Xd_0__inst_mult_20_11_q ;
wire Xd_0__inst_mult_19_10_q ;
wire Xd_0__inst_mult_19_11_q ;
wire Xd_0__inst_mult_18_10_q ;
wire Xd_0__inst_mult_18_11_q ;
wire Xd_0__inst_mult_17_10_q ;
wire Xd_0__inst_mult_17_11_q ;
wire Xd_0__inst_mult_16_10_q ;
wire Xd_0__inst_mult_16_11_q ;
wire Xd_0__inst_mult_15_10_q ;
wire Xd_0__inst_mult_15_11_q ;
wire Xd_0__inst_mult_14_10_q ;
wire Xd_0__inst_mult_14_11_q ;
wire Xd_0__inst_mult_13_10_q ;
wire Xd_0__inst_mult_13_11_q ;
wire Xd_0__inst_mult_12_10_q ;
wire Xd_0__inst_mult_12_11_q ;
wire Xd_0__inst_mult_11_10_q ;
wire Xd_0__inst_mult_11_11_q ;
wire Xd_0__inst_mult_10_10_q ;
wire Xd_0__inst_mult_10_11_q ;
wire Xd_0__inst_mult_9_10_q ;
wire Xd_0__inst_mult_9_11_q ;
wire Xd_0__inst_mult_8_10_q ;
wire Xd_0__inst_mult_8_11_q ;
wire Xd_0__inst_mult_7_10_q ;
wire Xd_0__inst_mult_7_11_q ;
wire Xd_0__inst_mult_6_10_q ;
wire Xd_0__inst_mult_6_11_q ;
wire Xd_0__inst_mult_5_10_q ;
wire Xd_0__inst_mult_5_11_q ;
wire Xd_0__inst_mult_4_10_q ;
wire Xd_0__inst_mult_4_11_q ;
wire Xd_0__inst_mult_3_10_q ;
wire Xd_0__inst_mult_3_11_q ;
wire Xd_0__inst_mult_2_10_q ;
wire Xd_0__inst_mult_2_11_q ;
wire Xd_0__inst_mult_1_10_q ;
wire Xd_0__inst_mult_1_11_q ;
wire Xd_0__inst_mult_0_10_q ;
wire Xd_0__inst_mult_0_11_q ;
wire Xd_0__inst_mult_31_12_q ;
wire Xd_0__inst_mult_31_13_q ;
wire Xd_0__inst_mult_31_14_q ;
wire Xd_0__inst_mult_31_15_q ;
wire Xd_0__inst_mult_30_12_q ;
wire Xd_0__inst_mult_30_13_q ;
wire Xd_0__inst_mult_30_14_q ;
wire Xd_0__inst_mult_30_15_q ;
wire Xd_0__inst_mult_29_12_q ;
wire Xd_0__inst_mult_29_13_q ;
wire Xd_0__inst_mult_29_14_q ;
wire Xd_0__inst_mult_29_15_q ;
wire Xd_0__inst_mult_28_12_q ;
wire Xd_0__inst_mult_28_13_q ;
wire Xd_0__inst_mult_28_14_q ;
wire Xd_0__inst_mult_28_15_q ;
wire Xd_0__inst_mult_27_12_q ;
wire Xd_0__inst_mult_27_13_q ;
wire Xd_0__inst_mult_27_14_q ;
wire Xd_0__inst_mult_27_15_q ;
wire Xd_0__inst_mult_26_12_q ;
wire Xd_0__inst_mult_26_13_q ;
wire Xd_0__inst_mult_26_14_q ;
wire Xd_0__inst_mult_26_15_q ;
wire Xd_0__inst_mult_25_12_q ;
wire Xd_0__inst_mult_25_13_q ;
wire Xd_0__inst_mult_25_14_q ;
wire Xd_0__inst_mult_25_15_q ;
wire Xd_0__inst_mult_24_12_q ;
wire Xd_0__inst_mult_24_13_q ;
wire Xd_0__inst_mult_24_14_q ;
wire Xd_0__inst_mult_24_15_q ;
wire Xd_0__inst_mult_23_12_q ;
wire Xd_0__inst_mult_23_13_q ;
wire Xd_0__inst_mult_23_14_q ;
wire Xd_0__inst_mult_23_15_q ;
wire Xd_0__inst_mult_22_12_q ;
wire Xd_0__inst_mult_22_13_q ;
wire Xd_0__inst_mult_22_14_q ;
wire Xd_0__inst_mult_22_15_q ;
wire Xd_0__inst_mult_21_12_q ;
wire Xd_0__inst_mult_21_13_q ;
wire Xd_0__inst_mult_21_14_q ;
wire Xd_0__inst_mult_21_15_q ;
wire Xd_0__inst_mult_20_12_q ;
wire Xd_0__inst_mult_20_13_q ;
wire Xd_0__inst_mult_20_14_q ;
wire Xd_0__inst_mult_20_15_q ;
wire Xd_0__inst_mult_19_12_q ;
wire Xd_0__inst_mult_19_13_q ;
wire Xd_0__inst_mult_19_14_q ;
wire Xd_0__inst_mult_19_15_q ;
wire Xd_0__inst_mult_18_12_q ;
wire Xd_0__inst_mult_18_13_q ;
wire Xd_0__inst_mult_18_14_q ;
wire Xd_0__inst_mult_18_15_q ;
wire Xd_0__inst_mult_17_12_q ;
wire Xd_0__inst_mult_17_13_q ;
wire Xd_0__inst_mult_17_14_q ;
wire Xd_0__inst_mult_17_15_q ;
wire Xd_0__inst_mult_16_12_q ;
wire Xd_0__inst_mult_16_13_q ;
wire Xd_0__inst_mult_16_14_q ;
wire Xd_0__inst_mult_16_15_q ;
wire Xd_0__inst_mult_15_12_q ;
wire Xd_0__inst_mult_15_13_q ;
wire Xd_0__inst_mult_15_14_q ;
wire Xd_0__inst_mult_15_15_q ;
wire Xd_0__inst_mult_14_12_q ;
wire Xd_0__inst_mult_14_13_q ;
wire Xd_0__inst_mult_14_14_q ;
wire Xd_0__inst_mult_14_15_q ;
wire Xd_0__inst_mult_13_12_q ;
wire Xd_0__inst_mult_13_13_q ;
wire Xd_0__inst_mult_13_14_q ;
wire Xd_0__inst_mult_13_15_q ;
wire Xd_0__inst_mult_12_12_q ;
wire Xd_0__inst_mult_12_13_q ;
wire Xd_0__inst_mult_12_14_q ;
wire Xd_0__inst_mult_12_15_q ;
wire Xd_0__inst_mult_11_12_q ;
wire Xd_0__inst_mult_11_13_q ;
wire Xd_0__inst_mult_11_14_q ;
wire Xd_0__inst_mult_11_15_q ;
wire Xd_0__inst_mult_10_12_q ;
wire Xd_0__inst_mult_10_13_q ;
wire Xd_0__inst_mult_10_14_q ;
wire Xd_0__inst_mult_10_15_q ;
wire Xd_0__inst_mult_9_12_q ;
wire Xd_0__inst_mult_9_13_q ;
wire Xd_0__inst_mult_9_14_q ;
wire Xd_0__inst_mult_9_15_q ;
wire Xd_0__inst_mult_8_12_q ;
wire Xd_0__inst_mult_8_13_q ;
wire Xd_0__inst_mult_8_14_q ;
wire Xd_0__inst_mult_8_15_q ;
wire Xd_0__inst_mult_7_12_q ;
wire Xd_0__inst_mult_7_13_q ;
wire Xd_0__inst_mult_7_14_q ;
wire Xd_0__inst_mult_7_15_q ;
wire Xd_0__inst_mult_6_12_q ;
wire Xd_0__inst_mult_6_13_q ;
wire Xd_0__inst_mult_6_14_q ;
wire Xd_0__inst_mult_6_15_q ;
wire Xd_0__inst_mult_5_12_q ;
wire Xd_0__inst_mult_5_13_q ;
wire Xd_0__inst_mult_5_14_q ;
wire Xd_0__inst_mult_5_15_q ;
wire Xd_0__inst_mult_4_12_q ;
wire Xd_0__inst_mult_4_13_q ;
wire Xd_0__inst_mult_4_14_q ;
wire Xd_0__inst_mult_4_15_q ;
wire Xd_0__inst_mult_3_12_q ;
wire Xd_0__inst_mult_3_13_q ;
wire Xd_0__inst_mult_3_14_q ;
wire Xd_0__inst_mult_3_15_q ;
wire Xd_0__inst_mult_2_12_q ;
wire Xd_0__inst_mult_2_13_q ;
wire Xd_0__inst_mult_2_14_q ;
wire Xd_0__inst_mult_2_15_q ;
wire Xd_0__inst_mult_1_12_q ;
wire Xd_0__inst_mult_1_13_q ;
wire Xd_0__inst_mult_1_14_q ;
wire Xd_0__inst_mult_1_15_q ;
wire Xd_0__inst_mult_0_12_q ;
wire Xd_0__inst_mult_0_13_q ;
wire Xd_0__inst_mult_0_14_q ;
wire Xd_0__inst_mult_0_15_q ;
wire Xd_0__inst_mult_31_16_q ;
wire Xd_0__inst_mult_31_17_q ;
wire Xd_0__inst_mult_30_16_q ;
wire Xd_0__inst_mult_30_17_q ;
wire Xd_0__inst_mult_29_16_q ;
wire Xd_0__inst_mult_29_17_q ;
wire Xd_0__inst_mult_28_16_q ;
wire Xd_0__inst_mult_28_17_q ;
wire Xd_0__inst_mult_27_16_q ;
wire Xd_0__inst_mult_27_17_q ;
wire Xd_0__inst_mult_26_16_q ;
wire Xd_0__inst_mult_26_17_q ;
wire Xd_0__inst_mult_25_16_q ;
wire Xd_0__inst_mult_25_17_q ;
wire Xd_0__inst_mult_24_16_q ;
wire Xd_0__inst_mult_24_17_q ;
wire Xd_0__inst_mult_23_16_q ;
wire Xd_0__inst_mult_23_17_q ;
wire Xd_0__inst_mult_22_16_q ;
wire Xd_0__inst_mult_22_17_q ;
wire Xd_0__inst_mult_21_16_q ;
wire Xd_0__inst_mult_21_17_q ;
wire Xd_0__inst_mult_20_16_q ;
wire Xd_0__inst_mult_20_17_q ;
wire Xd_0__inst_mult_19_16_q ;
wire Xd_0__inst_mult_19_17_q ;
wire Xd_0__inst_mult_18_16_q ;
wire Xd_0__inst_mult_18_17_q ;
wire Xd_0__inst_mult_17_16_q ;
wire Xd_0__inst_mult_17_17_q ;
wire Xd_0__inst_mult_16_16_q ;
wire Xd_0__inst_mult_16_17_q ;
wire Xd_0__inst_mult_15_16_q ;
wire Xd_0__inst_mult_15_17_q ;
wire Xd_0__inst_mult_14_16_q ;
wire Xd_0__inst_mult_14_17_q ;
wire Xd_0__inst_mult_13_16_q ;
wire Xd_0__inst_mult_13_17_q ;
wire Xd_0__inst_mult_12_16_q ;
wire Xd_0__inst_mult_12_17_q ;
wire Xd_0__inst_mult_11_16_q ;
wire Xd_0__inst_mult_11_17_q ;
wire Xd_0__inst_mult_10_16_q ;
wire Xd_0__inst_mult_10_17_q ;
wire Xd_0__inst_mult_9_16_q ;
wire Xd_0__inst_mult_9_17_q ;
wire Xd_0__inst_mult_8_16_q ;
wire Xd_0__inst_mult_8_17_q ;
wire Xd_0__inst_mult_7_16_q ;
wire Xd_0__inst_mult_7_17_q ;
wire Xd_0__inst_mult_6_16_q ;
wire Xd_0__inst_mult_6_17_q ;
wire Xd_0__inst_mult_5_16_q ;
wire Xd_0__inst_mult_5_17_q ;
wire Xd_0__inst_mult_4_16_q ;
wire Xd_0__inst_mult_4_17_q ;
wire Xd_0__inst_mult_3_16_q ;
wire Xd_0__inst_mult_3_17_q ;
wire Xd_0__inst_mult_2_16_q ;
wire Xd_0__inst_mult_2_17_q ;
wire Xd_0__inst_mult_1_16_q ;
wire Xd_0__inst_mult_1_17_q ;
wire Xd_0__inst_mult_0_16_q ;
wire Xd_0__inst_mult_0_17_q ;
wire Xd_0__inst_mult_31_18_q ;
wire Xd_0__inst_mult_31_19_q ;
wire Xd_0__inst_mult_30_18_q ;
wire Xd_0__inst_mult_30_19_q ;
wire Xd_0__inst_mult_29_18_q ;
wire Xd_0__inst_mult_29_19_q ;
wire Xd_0__inst_mult_28_18_q ;
wire Xd_0__inst_mult_28_19_q ;
wire Xd_0__inst_mult_27_18_q ;
wire Xd_0__inst_mult_27_19_q ;
wire Xd_0__inst_mult_26_18_q ;
wire Xd_0__inst_mult_26_19_q ;
wire Xd_0__inst_mult_25_18_q ;
wire Xd_0__inst_mult_25_19_q ;
wire Xd_0__inst_mult_24_18_q ;
wire Xd_0__inst_mult_24_19_q ;
wire Xd_0__inst_mult_23_18_q ;
wire Xd_0__inst_mult_23_19_q ;
wire Xd_0__inst_mult_22_18_q ;
wire Xd_0__inst_mult_22_19_q ;
wire Xd_0__inst_mult_21_18_q ;
wire Xd_0__inst_mult_21_19_q ;
wire Xd_0__inst_mult_20_18_q ;
wire Xd_0__inst_mult_20_19_q ;
wire Xd_0__inst_mult_19_18_q ;
wire Xd_0__inst_mult_19_19_q ;
wire Xd_0__inst_mult_18_18_q ;
wire Xd_0__inst_mult_18_19_q ;
wire Xd_0__inst_mult_17_18_q ;
wire Xd_0__inst_mult_17_19_q ;
wire Xd_0__inst_mult_16_18_q ;
wire Xd_0__inst_mult_16_19_q ;
wire Xd_0__inst_mult_15_18_q ;
wire Xd_0__inst_mult_15_19_q ;
wire Xd_0__inst_mult_14_18_q ;
wire Xd_0__inst_mult_14_19_q ;
wire Xd_0__inst_mult_13_18_q ;
wire Xd_0__inst_mult_13_19_q ;
wire Xd_0__inst_mult_12_18_q ;
wire Xd_0__inst_mult_12_19_q ;
wire Xd_0__inst_mult_11_18_q ;
wire Xd_0__inst_mult_11_19_q ;
wire Xd_0__inst_mult_10_18_q ;
wire Xd_0__inst_mult_10_19_q ;
wire Xd_0__inst_mult_9_18_q ;
wire Xd_0__inst_mult_9_19_q ;
wire Xd_0__inst_mult_8_18_q ;
wire Xd_0__inst_mult_8_19_q ;
wire Xd_0__inst_mult_7_18_q ;
wire Xd_0__inst_mult_7_19_q ;
wire Xd_0__inst_mult_6_18_q ;
wire Xd_0__inst_mult_6_19_q ;
wire Xd_0__inst_mult_5_18_q ;
wire Xd_0__inst_mult_5_19_q ;
wire Xd_0__inst_mult_4_18_q ;
wire Xd_0__inst_mult_4_19_q ;
wire Xd_0__inst_mult_3_18_q ;
wire Xd_0__inst_mult_3_19_q ;
wire Xd_0__inst_mult_2_18_q ;
wire Xd_0__inst_mult_2_19_q ;
wire Xd_0__inst_mult_1_18_q ;
wire Xd_0__inst_mult_1_19_q ;
wire Xd_0__inst_mult_0_18_q ;
wire Xd_0__inst_mult_0_19_q ;
wire Xd_0__inst_mult_31_20_q ;
wire Xd_0__inst_mult_31_21_q ;
wire Xd_0__inst_mult_30_20_q ;
wire Xd_0__inst_mult_30_21_q ;
wire Xd_0__inst_mult_29_20_q ;
wire Xd_0__inst_mult_29_21_q ;
wire Xd_0__inst_mult_28_20_q ;
wire Xd_0__inst_mult_28_21_q ;
wire Xd_0__inst_mult_27_20_q ;
wire Xd_0__inst_mult_27_21_q ;
wire Xd_0__inst_mult_26_20_q ;
wire Xd_0__inst_mult_26_21_q ;
wire Xd_0__inst_mult_25_20_q ;
wire Xd_0__inst_mult_25_21_q ;
wire Xd_0__inst_mult_24_20_q ;
wire Xd_0__inst_mult_24_21_q ;
wire Xd_0__inst_mult_23_20_q ;
wire Xd_0__inst_mult_23_21_q ;
wire Xd_0__inst_mult_22_20_q ;
wire Xd_0__inst_mult_22_21_q ;
wire Xd_0__inst_mult_21_20_q ;
wire Xd_0__inst_mult_21_21_q ;
wire Xd_0__inst_mult_20_20_q ;
wire Xd_0__inst_mult_20_21_q ;
wire Xd_0__inst_mult_19_20_q ;
wire Xd_0__inst_mult_19_21_q ;
wire Xd_0__inst_mult_18_20_q ;
wire Xd_0__inst_mult_18_21_q ;
wire Xd_0__inst_mult_17_20_q ;
wire Xd_0__inst_mult_17_21_q ;
wire Xd_0__inst_mult_16_20_q ;
wire Xd_0__inst_mult_16_21_q ;
wire Xd_0__inst_mult_15_20_q ;
wire Xd_0__inst_mult_15_21_q ;
wire Xd_0__inst_mult_14_20_q ;
wire Xd_0__inst_mult_14_21_q ;
wire Xd_0__inst_mult_13_20_q ;
wire Xd_0__inst_mult_13_21_q ;
wire Xd_0__inst_mult_12_20_q ;
wire Xd_0__inst_mult_12_21_q ;
wire Xd_0__inst_mult_11_20_q ;
wire Xd_0__inst_mult_11_21_q ;
wire Xd_0__inst_mult_10_20_q ;
wire Xd_0__inst_mult_10_21_q ;
wire Xd_0__inst_mult_9_20_q ;
wire Xd_0__inst_mult_9_21_q ;
wire Xd_0__inst_mult_8_20_q ;
wire Xd_0__inst_mult_8_21_q ;
wire Xd_0__inst_mult_7_20_q ;
wire Xd_0__inst_mult_7_21_q ;
wire Xd_0__inst_mult_6_20_q ;
wire Xd_0__inst_mult_6_21_q ;
wire Xd_0__inst_mult_5_20_q ;
wire Xd_0__inst_mult_5_21_q ;
wire Xd_0__inst_mult_4_20_q ;
wire Xd_0__inst_mult_4_21_q ;
wire Xd_0__inst_mult_3_20_q ;
wire Xd_0__inst_mult_3_21_q ;
wire Xd_0__inst_mult_2_20_q ;
wire Xd_0__inst_mult_2_21_q ;
wire Xd_0__inst_mult_1_20_q ;
wire Xd_0__inst_mult_1_21_q ;
wire Xd_0__inst_mult_0_20_q ;
wire Xd_0__inst_mult_0_21_q ;
wire [0:31] Xd_0__inst_sign1 ;
wire [0:31] Xd_0__inst_sign ;
wire [0:15] Xd_0__inst_r_sign ;
wire [19:0] Xd_0__inst_inst_inst_inst_dout ;


fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__14__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__16__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__17__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_inst_inst_first_level_1__18__q ),
	.datab(!Xd_0__inst_inst_inst_first_level_0__18__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_inst_inst_first_level_1__18__q ),
	.datab(!Xd_0__inst_inst_inst_first_level_0__18__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_96_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__0__q ),
	.datad(!Xd_0__inst_inst_first_level_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__1__q ),
	.datad(!Xd_0__inst_inst_first_level_2__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_6_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__2__q ),
	.datad(!Xd_0__inst_inst_first_level_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_11_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__3__q ),
	.datad(!Xd_0__inst_inst_first_level_2__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_16_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__4__q ),
	.datad(!Xd_0__inst_inst_first_level_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__5__q ),
	.datad(!Xd_0__inst_inst_first_level_2__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_26_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__6__q ),
	.datad(!Xd_0__inst_inst_first_level_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_31_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__7__q ),
	.datad(!Xd_0__inst_inst_first_level_2__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_36_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__8__q ),
	.datad(!Xd_0__inst_inst_first_level_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__9__q ),
	.datad(!Xd_0__inst_inst_first_level_2__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_46_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__10__q ),
	.datad(!Xd_0__inst_inst_first_level_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_51_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__11__q ),
	.datad(!Xd_0__inst_inst_first_level_2__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_56_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__12__q ),
	.datad(!Xd_0__inst_inst_first_level_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__13__q ),
	.datad(!Xd_0__inst_inst_first_level_2__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_66_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__14__q ),
	.datad(!Xd_0__inst_inst_first_level_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_71_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__14__q ),
	.datad(!Xd_0__inst_inst_first_level_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__15__q ),
	.datad(!Xd_0__inst_inst_first_level_2__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_76_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__16__q ),
	.datad(!Xd_0__inst_inst_first_level_2__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_81_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__16__q ),
	.datad(!Xd_0__inst_inst_first_level_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__17__q ),
	.datad(!Xd_0__inst_inst_first_level_2__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_86_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__17__q ),
	.datad(!Xd_0__inst_inst_first_level_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__17__q ),
	.datad(!Xd_0__inst_inst_first_level_2__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_91_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__17__q ),
	.datad(!Xd_0__inst_inst_first_level_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_91_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_23 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[101]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_23_sumout ),
	.cout(Xd_0__inst_mult_12_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_23 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[109]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_23_sumout ),
	.cout(Xd_0__inst_mult_13_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__0__q ),
	.datad(!Xd_0__inst_r_sum2_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_1_sumout ),
	.cout(Xd_0__inst_inst_add_3_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__0__q ),
	.datad(!Xd_0__inst_r_sum2_4__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_1_sumout ),
	.cout(Xd_0__inst_inst_add_2_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__0__q ),
	.datad(!Xd_0__inst_r_sum2_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_1_sumout ),
	.cout(Xd_0__inst_inst_add_1_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__0__q ),
	.datad(!Xd_0__inst_r_sum2_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__1__q ),
	.datad(!Xd_0__inst_r_sum2_6__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_6_sumout ),
	.cout(Xd_0__inst_inst_add_3_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__1__q ),
	.datad(!Xd_0__inst_r_sum2_4__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_6_sumout ),
	.cout(Xd_0__inst_inst_add_2_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__1__q ),
	.datad(!Xd_0__inst_r_sum2_2__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_6_sumout ),
	.cout(Xd_0__inst_inst_add_1_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__1__q ),
	.datad(!Xd_0__inst_r_sum2_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__2__q ),
	.datad(!Xd_0__inst_r_sum2_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_11_sumout ),
	.cout(Xd_0__inst_inst_add_3_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__2__q ),
	.datad(!Xd_0__inst_r_sum2_4__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_11_sumout ),
	.cout(Xd_0__inst_inst_add_2_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__2__q ),
	.datad(!Xd_0__inst_r_sum2_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_11_sumout ),
	.cout(Xd_0__inst_inst_add_1_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__2__q ),
	.datad(!Xd_0__inst_r_sum2_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__3__q ),
	.datad(!Xd_0__inst_r_sum2_6__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_16_sumout ),
	.cout(Xd_0__inst_inst_add_3_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__3__q ),
	.datad(!Xd_0__inst_r_sum2_4__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_16_sumout ),
	.cout(Xd_0__inst_inst_add_2_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__3__q ),
	.datad(!Xd_0__inst_r_sum2_2__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_16_sumout ),
	.cout(Xd_0__inst_inst_add_1_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__3__q ),
	.datad(!Xd_0__inst_r_sum2_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__4__q ),
	.datad(!Xd_0__inst_r_sum2_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_21_sumout ),
	.cout(Xd_0__inst_inst_add_3_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__4__q ),
	.datad(!Xd_0__inst_r_sum2_4__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_21_sumout ),
	.cout(Xd_0__inst_inst_add_2_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__4__q ),
	.datad(!Xd_0__inst_r_sum2_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_21_sumout ),
	.cout(Xd_0__inst_inst_add_1_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__4__q ),
	.datad(!Xd_0__inst_r_sum2_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__5__q ),
	.datad(!Xd_0__inst_r_sum2_6__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_26_sumout ),
	.cout(Xd_0__inst_inst_add_3_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__5__q ),
	.datad(!Xd_0__inst_r_sum2_4__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_26_sumout ),
	.cout(Xd_0__inst_inst_add_2_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__5__q ),
	.datad(!Xd_0__inst_r_sum2_2__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_26_sumout ),
	.cout(Xd_0__inst_inst_add_1_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__5__q ),
	.datad(!Xd_0__inst_r_sum2_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__6__q ),
	.datad(!Xd_0__inst_r_sum2_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_31_sumout ),
	.cout(Xd_0__inst_inst_add_3_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__6__q ),
	.datad(!Xd_0__inst_r_sum2_4__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_31_sumout ),
	.cout(Xd_0__inst_inst_add_2_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__6__q ),
	.datad(!Xd_0__inst_r_sum2_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_31_sumout ),
	.cout(Xd_0__inst_inst_add_1_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__6__q ),
	.datad(!Xd_0__inst_r_sum2_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__7__q ),
	.datad(!Xd_0__inst_r_sum2_6__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_36_sumout ),
	.cout(Xd_0__inst_inst_add_3_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__7__q ),
	.datad(!Xd_0__inst_r_sum2_4__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_36_sumout ),
	.cout(Xd_0__inst_inst_add_2_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__7__q ),
	.datad(!Xd_0__inst_r_sum2_2__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_36_sumout ),
	.cout(Xd_0__inst_inst_add_1_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__7__q ),
	.datad(!Xd_0__inst_r_sum2_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__8__q ),
	.datad(!Xd_0__inst_r_sum2_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_41_sumout ),
	.cout(Xd_0__inst_inst_add_3_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__8__q ),
	.datad(!Xd_0__inst_r_sum2_4__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_41_sumout ),
	.cout(Xd_0__inst_inst_add_2_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__8__q ),
	.datad(!Xd_0__inst_r_sum2_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_41_sumout ),
	.cout(Xd_0__inst_inst_add_1_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__8__q ),
	.datad(!Xd_0__inst_r_sum2_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__9__q ),
	.datad(!Xd_0__inst_r_sum2_6__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_46_sumout ),
	.cout(Xd_0__inst_inst_add_3_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__9__q ),
	.datad(!Xd_0__inst_r_sum2_4__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_46_sumout ),
	.cout(Xd_0__inst_inst_add_2_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__9__q ),
	.datad(!Xd_0__inst_r_sum2_2__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_46_sumout ),
	.cout(Xd_0__inst_inst_add_1_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__9__q ),
	.datad(!Xd_0__inst_r_sum2_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__10__q ),
	.datad(!Xd_0__inst_r_sum2_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_51_sumout ),
	.cout(Xd_0__inst_inst_add_3_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__10__q ),
	.datad(!Xd_0__inst_r_sum2_4__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_51_sumout ),
	.cout(Xd_0__inst_inst_add_2_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__10__q ),
	.datad(!Xd_0__inst_r_sum2_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_51_sumout ),
	.cout(Xd_0__inst_inst_add_1_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__10__q ),
	.datad(!Xd_0__inst_r_sum2_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__11__q ),
	.datad(!Xd_0__inst_r_sum2_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_56_sumout ),
	.cout(Xd_0__inst_inst_add_3_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__11__q ),
	.datad(!Xd_0__inst_r_sum2_4__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_56_sumout ),
	.cout(Xd_0__inst_inst_add_2_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__11__q ),
	.datad(!Xd_0__inst_r_sum2_2__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_56_sumout ),
	.cout(Xd_0__inst_inst_add_1_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__11__q ),
	.datad(!Xd_0__inst_r_sum2_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__12__q ),
	.datad(!Xd_0__inst_r_sum2_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_61_sumout ),
	.cout(Xd_0__inst_inst_add_3_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__12__q ),
	.datad(!Xd_0__inst_r_sum2_4__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_61_sumout ),
	.cout(Xd_0__inst_inst_add_2_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__12__q ),
	.datad(!Xd_0__inst_r_sum2_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_61_sumout ),
	.cout(Xd_0__inst_inst_add_1_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__12__q ),
	.datad(!Xd_0__inst_r_sum2_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__13__q ),
	.datad(!Xd_0__inst_r_sum2_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_66_sumout ),
	.cout(Xd_0__inst_inst_add_3_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__13__q ),
	.datad(!Xd_0__inst_r_sum2_4__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_66_sumout ),
	.cout(Xd_0__inst_inst_add_2_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__13__q ),
	.datad(!Xd_0__inst_r_sum2_2__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_66_sumout ),
	.cout(Xd_0__inst_inst_add_1_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__13__q ),
	.datad(!Xd_0__inst_r_sum2_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__14__q ),
	.datad(!Xd_0__inst_r_sum2_6__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_71_sumout ),
	.cout(Xd_0__inst_inst_add_3_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__14__q ),
	.datad(!Xd_0__inst_r_sum2_4__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_71_sumout ),
	.cout(Xd_0__inst_inst_add_2_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__14__q ),
	.datad(!Xd_0__inst_r_sum2_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_71_sumout ),
	.cout(Xd_0__inst_inst_add_1_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__14__q ),
	.datad(!Xd_0__inst_r_sum2_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__15__q ),
	.datad(!Xd_0__inst_r_sum2_6__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_76_sumout ),
	.cout(Xd_0__inst_inst_add_3_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__15__q ),
	.datad(!Xd_0__inst_r_sum2_4__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_76_sumout ),
	.cout(Xd_0__inst_inst_add_2_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__15__q ),
	.datad(!Xd_0__inst_r_sum2_2__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_76_sumout ),
	.cout(Xd_0__inst_inst_add_1_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__15__q ),
	.datad(!Xd_0__inst_r_sum2_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_7__16__q ),
	.datab(!Xd_0__inst_r_sum2_6__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_81_sumout ),
	.cout(Xd_0__inst_inst_add_3_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_5__16__q ),
	.datab(!Xd_0__inst_r_sum2_4__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_81_sumout ),
	.cout(Xd_0__inst_inst_add_2_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_3__16__q ),
	.datab(!Xd_0__inst_r_sum2_2__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_81_sumout ),
	.cout(Xd_0__inst_inst_add_1_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_1__16__q ),
	.datab(!Xd_0__inst_r_sum2_0__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_7__16__q ),
	.datab(!Xd_0__inst_r_sum2_6__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_86_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_5__16__q ),
	.datab(!Xd_0__inst_r_sum2_4__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_86_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_3__16__q ),
	.datab(!Xd_0__inst_r_sum2_2__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_86_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_1__16__q ),
	.datab(!Xd_0__inst_r_sum2_0__16__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_86_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_23 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_23_sumout ),
	.cout(Xd_0__inst_mult_11_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_23 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[181]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_23_sumout ),
	.cout(Xd_0__inst_mult_22_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_23 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[197]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_23_sumout ),
	.cout(Xd_0__inst_mult_24_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_23 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[213]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_23_sumout ),
	.cout(Xd_0__inst_mult_26_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_14__0__q ),
	.datad(!Xd_0__inst_r_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_12__0__q ),
	.datad(!Xd_0__inst_r_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_23 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[85]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_23_sumout ),
	.cout(Xd_0__inst_mult_10_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_10__0__q ),
	.datad(!Xd_0__inst_r_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_8__0__q ),
	.datad(!Xd_0__inst_r_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_23 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[173]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_23_sumout ),
	.cout(Xd_0__inst_mult_21_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_6__0__q ),
	.datad(!Xd_0__inst_r_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_4__0__q ),
	.datad(!Xd_0__inst_r_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_23 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[117]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_23_sumout ),
	.cout(Xd_0__inst_mult_14_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_2__0__q ),
	.datad(!Xd_0__inst_r_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_0__0__q ),
	.datad(!Xd_0__inst_r_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_87_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_23 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[205]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_23_sumout ),
	.cout(Xd_0__inst_mult_25_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__1__q ),
	.datab(!Xd_0__inst_r_sum1_14__1__q ),
	.datac(!Xd_0__inst_r_sum1_14__0__q ),
	.datad(!Xd_0__inst_r_sum1_15__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__1__q ),
	.datab(!Xd_0__inst_r_sum1_12__1__q ),
	.datac(!Xd_0__inst_r_sum1_12__0__q ),
	.datad(!Xd_0__inst_r_sum1_13__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__1__q ),
	.datab(!Xd_0__inst_r_sum1_10__1__q ),
	.datac(!Xd_0__inst_r_sum1_10__0__q ),
	.datad(!Xd_0__inst_r_sum1_11__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__1__q ),
	.datab(!Xd_0__inst_r_sum1_8__1__q ),
	.datac(!Xd_0__inst_r_sum1_8__0__q ),
	.datad(!Xd_0__inst_r_sum1_9__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__1__q ),
	.datab(!Xd_0__inst_r_sum1_6__1__q ),
	.datac(!Xd_0__inst_r_sum1_6__0__q ),
	.datad(!Xd_0__inst_r_sum1_7__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__1__q ),
	.datab(!Xd_0__inst_r_sum1_4__1__q ),
	.datac(!Xd_0__inst_r_sum1_4__0__q ),
	.datad(!Xd_0__inst_r_sum1_5__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__1__q ),
	.datab(!Xd_0__inst_r_sum1_2__1__q ),
	.datac(!Xd_0__inst_r_sum1_2__0__q ),
	.datad(!Xd_0__inst_r_sum1_3__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__1__q ),
	.datab(!Xd_0__inst_r_sum1_0__1__q ),
	.datac(!Xd_0__inst_r_sum1_0__0__q ),
	.datad(!Xd_0__inst_r_sum1_1__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__1__q ),
	.datab(!Xd_0__inst_r_sum1_14__1__q ),
	.datac(!Xd_0__inst_r_sum1_15__2__q ),
	.datad(!Xd_0__inst_r_sum1_14__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__1__q ),
	.datab(!Xd_0__inst_r_sum1_12__1__q ),
	.datac(!Xd_0__inst_r_sum1_13__2__q ),
	.datad(!Xd_0__inst_r_sum1_12__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__1__q ),
	.datab(!Xd_0__inst_r_sum1_10__1__q ),
	.datac(!Xd_0__inst_r_sum1_11__2__q ),
	.datad(!Xd_0__inst_r_sum1_10__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__1__q ),
	.datab(!Xd_0__inst_r_sum1_8__1__q ),
	.datac(!Xd_0__inst_r_sum1_9__2__q ),
	.datad(!Xd_0__inst_r_sum1_8__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__1__q ),
	.datab(!Xd_0__inst_r_sum1_6__1__q ),
	.datac(!Xd_0__inst_r_sum1_7__2__q ),
	.datad(!Xd_0__inst_r_sum1_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__1__q ),
	.datab(!Xd_0__inst_r_sum1_4__1__q ),
	.datac(!Xd_0__inst_r_sum1_5__2__q ),
	.datad(!Xd_0__inst_r_sum1_4__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__1__q ),
	.datab(!Xd_0__inst_r_sum1_2__1__q ),
	.datac(!Xd_0__inst_r_sum1_3__2__q ),
	.datad(!Xd_0__inst_r_sum1_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__1__q ),
	.datab(!Xd_0__inst_r_sum1_0__1__q ),
	.datac(!Xd_0__inst_r_sum1_1__2__q ),
	.datad(!Xd_0__inst_r_sum1_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__3__q ),
	.datab(!Xd_0__inst_r_sum1_14__3__q ),
	.datac(!Xd_0__inst_r_sum1_14__2__q ),
	.datad(!Xd_0__inst_r_sum1_15__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__3__q ),
	.datab(!Xd_0__inst_r_sum1_12__3__q ),
	.datac(!Xd_0__inst_r_sum1_12__2__q ),
	.datad(!Xd_0__inst_r_sum1_13__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__3__q ),
	.datab(!Xd_0__inst_r_sum1_10__3__q ),
	.datac(!Xd_0__inst_r_sum1_10__2__q ),
	.datad(!Xd_0__inst_r_sum1_11__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__3__q ),
	.datab(!Xd_0__inst_r_sum1_8__3__q ),
	.datac(!Xd_0__inst_r_sum1_8__2__q ),
	.datad(!Xd_0__inst_r_sum1_9__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__3__q ),
	.datab(!Xd_0__inst_r_sum1_6__3__q ),
	.datac(!Xd_0__inst_r_sum1_6__2__q ),
	.datad(!Xd_0__inst_r_sum1_7__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__3__q ),
	.datab(!Xd_0__inst_r_sum1_4__3__q ),
	.datac(!Xd_0__inst_r_sum1_4__2__q ),
	.datad(!Xd_0__inst_r_sum1_5__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__3__q ),
	.datab(!Xd_0__inst_r_sum1_2__3__q ),
	.datac(!Xd_0__inst_r_sum1_2__2__q ),
	.datad(!Xd_0__inst_r_sum1_3__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__3__q ),
	.datab(!Xd_0__inst_r_sum1_0__3__q ),
	.datac(!Xd_0__inst_r_sum1_0__2__q ),
	.datad(!Xd_0__inst_r_sum1_1__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__3__q ),
	.datab(!Xd_0__inst_r_sum1_14__3__q ),
	.datac(!Xd_0__inst_r_sum1_15__4__q ),
	.datad(!Xd_0__inst_r_sum1_14__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__3__q ),
	.datab(!Xd_0__inst_r_sum1_12__3__q ),
	.datac(!Xd_0__inst_r_sum1_13__4__q ),
	.datad(!Xd_0__inst_r_sum1_12__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__3__q ),
	.datab(!Xd_0__inst_r_sum1_10__3__q ),
	.datac(!Xd_0__inst_r_sum1_11__4__q ),
	.datad(!Xd_0__inst_r_sum1_10__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__3__q ),
	.datab(!Xd_0__inst_r_sum1_8__3__q ),
	.datac(!Xd_0__inst_r_sum1_9__4__q ),
	.datad(!Xd_0__inst_r_sum1_8__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__3__q ),
	.datab(!Xd_0__inst_r_sum1_6__3__q ),
	.datac(!Xd_0__inst_r_sum1_7__4__q ),
	.datad(!Xd_0__inst_r_sum1_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__3__q ),
	.datab(!Xd_0__inst_r_sum1_4__3__q ),
	.datac(!Xd_0__inst_r_sum1_5__4__q ),
	.datad(!Xd_0__inst_r_sum1_4__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__3__q ),
	.datab(!Xd_0__inst_r_sum1_2__3__q ),
	.datac(!Xd_0__inst_r_sum1_3__4__q ),
	.datad(!Xd_0__inst_r_sum1_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__3__q ),
	.datab(!Xd_0__inst_r_sum1_0__3__q ),
	.datac(!Xd_0__inst_r_sum1_1__4__q ),
	.datad(!Xd_0__inst_r_sum1_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__5__q ),
	.datab(!Xd_0__inst_r_sum1_14__5__q ),
	.datac(!Xd_0__inst_r_sum1_14__4__q ),
	.datad(!Xd_0__inst_r_sum1_15__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__5__q ),
	.datab(!Xd_0__inst_r_sum1_12__5__q ),
	.datac(!Xd_0__inst_r_sum1_12__4__q ),
	.datad(!Xd_0__inst_r_sum1_13__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__5__q ),
	.datab(!Xd_0__inst_r_sum1_10__5__q ),
	.datac(!Xd_0__inst_r_sum1_10__4__q ),
	.datad(!Xd_0__inst_r_sum1_11__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__5__q ),
	.datab(!Xd_0__inst_r_sum1_8__5__q ),
	.datac(!Xd_0__inst_r_sum1_8__4__q ),
	.datad(!Xd_0__inst_r_sum1_9__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__5__q ),
	.datab(!Xd_0__inst_r_sum1_6__5__q ),
	.datac(!Xd_0__inst_r_sum1_6__4__q ),
	.datad(!Xd_0__inst_r_sum1_7__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__5__q ),
	.datab(!Xd_0__inst_r_sum1_4__5__q ),
	.datac(!Xd_0__inst_r_sum1_4__4__q ),
	.datad(!Xd_0__inst_r_sum1_5__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__5__q ),
	.datab(!Xd_0__inst_r_sum1_2__5__q ),
	.datac(!Xd_0__inst_r_sum1_2__4__q ),
	.datad(!Xd_0__inst_r_sum1_3__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__5__q ),
	.datab(!Xd_0__inst_r_sum1_0__5__q ),
	.datac(!Xd_0__inst_r_sum1_0__4__q ),
	.datad(!Xd_0__inst_r_sum1_1__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__5__q ),
	.datab(!Xd_0__inst_r_sum1_14__5__q ),
	.datac(!Xd_0__inst_r_sum1_15__6__q ),
	.datad(!Xd_0__inst_r_sum1_14__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__5__q ),
	.datab(!Xd_0__inst_r_sum1_12__5__q ),
	.datac(!Xd_0__inst_r_sum1_13__6__q ),
	.datad(!Xd_0__inst_r_sum1_12__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__5__q ),
	.datab(!Xd_0__inst_r_sum1_10__5__q ),
	.datac(!Xd_0__inst_r_sum1_11__6__q ),
	.datad(!Xd_0__inst_r_sum1_10__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__5__q ),
	.datab(!Xd_0__inst_r_sum1_8__5__q ),
	.datac(!Xd_0__inst_r_sum1_9__6__q ),
	.datad(!Xd_0__inst_r_sum1_8__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__5__q ),
	.datab(!Xd_0__inst_r_sum1_6__5__q ),
	.datac(!Xd_0__inst_r_sum1_7__6__q ),
	.datad(!Xd_0__inst_r_sum1_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__5__q ),
	.datab(!Xd_0__inst_r_sum1_4__5__q ),
	.datac(!Xd_0__inst_r_sum1_5__6__q ),
	.datad(!Xd_0__inst_r_sum1_4__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__5__q ),
	.datab(!Xd_0__inst_r_sum1_2__5__q ),
	.datac(!Xd_0__inst_r_sum1_3__6__q ),
	.datad(!Xd_0__inst_r_sum1_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__5__q ),
	.datab(!Xd_0__inst_r_sum1_0__5__q ),
	.datac(!Xd_0__inst_r_sum1_1__6__q ),
	.datad(!Xd_0__inst_r_sum1_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__7__q ),
	.datab(!Xd_0__inst_r_sum1_14__7__q ),
	.datac(!Xd_0__inst_r_sum1_14__6__q ),
	.datad(!Xd_0__inst_r_sum1_15__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__7__q ),
	.datab(!Xd_0__inst_r_sum1_12__7__q ),
	.datac(!Xd_0__inst_r_sum1_12__6__q ),
	.datad(!Xd_0__inst_r_sum1_13__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__7__q ),
	.datab(!Xd_0__inst_r_sum1_10__7__q ),
	.datac(!Xd_0__inst_r_sum1_10__6__q ),
	.datad(!Xd_0__inst_r_sum1_11__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__7__q ),
	.datab(!Xd_0__inst_r_sum1_8__7__q ),
	.datac(!Xd_0__inst_r_sum1_8__6__q ),
	.datad(!Xd_0__inst_r_sum1_9__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__7__q ),
	.datab(!Xd_0__inst_r_sum1_6__7__q ),
	.datac(!Xd_0__inst_r_sum1_6__6__q ),
	.datad(!Xd_0__inst_r_sum1_7__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__7__q ),
	.datab(!Xd_0__inst_r_sum1_4__7__q ),
	.datac(!Xd_0__inst_r_sum1_4__6__q ),
	.datad(!Xd_0__inst_r_sum1_5__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__7__q ),
	.datab(!Xd_0__inst_r_sum1_2__7__q ),
	.datac(!Xd_0__inst_r_sum1_2__6__q ),
	.datad(!Xd_0__inst_r_sum1_3__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__7__q ),
	.datab(!Xd_0__inst_r_sum1_0__7__q ),
	.datac(!Xd_0__inst_r_sum1_0__6__q ),
	.datad(!Xd_0__inst_r_sum1_1__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__7__q ),
	.datab(!Xd_0__inst_r_sum1_14__7__q ),
	.datac(!Xd_0__inst_r_sum1_15__8__q ),
	.datad(!Xd_0__inst_r_sum1_14__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__7__q ),
	.datab(!Xd_0__inst_r_sum1_12__7__q ),
	.datac(!Xd_0__inst_r_sum1_13__8__q ),
	.datad(!Xd_0__inst_r_sum1_12__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__7__q ),
	.datab(!Xd_0__inst_r_sum1_10__7__q ),
	.datac(!Xd_0__inst_r_sum1_11__8__q ),
	.datad(!Xd_0__inst_r_sum1_10__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__7__q ),
	.datab(!Xd_0__inst_r_sum1_8__7__q ),
	.datac(!Xd_0__inst_r_sum1_9__8__q ),
	.datad(!Xd_0__inst_r_sum1_8__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__7__q ),
	.datab(!Xd_0__inst_r_sum1_6__7__q ),
	.datac(!Xd_0__inst_r_sum1_7__8__q ),
	.datad(!Xd_0__inst_r_sum1_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__7__q ),
	.datab(!Xd_0__inst_r_sum1_4__7__q ),
	.datac(!Xd_0__inst_r_sum1_5__8__q ),
	.datad(!Xd_0__inst_r_sum1_4__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__7__q ),
	.datab(!Xd_0__inst_r_sum1_2__7__q ),
	.datac(!Xd_0__inst_r_sum1_3__8__q ),
	.datad(!Xd_0__inst_r_sum1_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__7__q ),
	.datab(!Xd_0__inst_r_sum1_0__7__q ),
	.datac(!Xd_0__inst_r_sum1_1__8__q ),
	.datad(!Xd_0__inst_r_sum1_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__9__q ),
	.datab(!Xd_0__inst_r_sum1_14__9__q ),
	.datac(!Xd_0__inst_r_sum1_14__8__q ),
	.datad(!Xd_0__inst_r_sum1_15__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__9__q ),
	.datab(!Xd_0__inst_r_sum1_12__9__q ),
	.datac(!Xd_0__inst_r_sum1_12__8__q ),
	.datad(!Xd_0__inst_r_sum1_13__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__9__q ),
	.datab(!Xd_0__inst_r_sum1_10__9__q ),
	.datac(!Xd_0__inst_r_sum1_10__8__q ),
	.datad(!Xd_0__inst_r_sum1_11__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__9__q ),
	.datab(!Xd_0__inst_r_sum1_8__9__q ),
	.datac(!Xd_0__inst_r_sum1_8__8__q ),
	.datad(!Xd_0__inst_r_sum1_9__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__9__q ),
	.datab(!Xd_0__inst_r_sum1_6__9__q ),
	.datac(!Xd_0__inst_r_sum1_6__8__q ),
	.datad(!Xd_0__inst_r_sum1_7__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__9__q ),
	.datab(!Xd_0__inst_r_sum1_4__9__q ),
	.datac(!Xd_0__inst_r_sum1_4__8__q ),
	.datad(!Xd_0__inst_r_sum1_5__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__9__q ),
	.datab(!Xd_0__inst_r_sum1_2__9__q ),
	.datac(!Xd_0__inst_r_sum1_2__8__q ),
	.datad(!Xd_0__inst_r_sum1_3__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__9__q ),
	.datab(!Xd_0__inst_r_sum1_0__9__q ),
	.datac(!Xd_0__inst_r_sum1_0__8__q ),
	.datad(!Xd_0__inst_r_sum1_1__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__9__q ),
	.datab(!Xd_0__inst_r_sum1_14__9__q ),
	.datac(!Xd_0__inst_r_sum1_15__10__q ),
	.datad(!Xd_0__inst_r_sum1_14__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__9__q ),
	.datab(!Xd_0__inst_r_sum1_12__9__q ),
	.datac(!Xd_0__inst_r_sum1_13__10__q ),
	.datad(!Xd_0__inst_r_sum1_12__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__9__q ),
	.datab(!Xd_0__inst_r_sum1_10__9__q ),
	.datac(!Xd_0__inst_r_sum1_11__10__q ),
	.datad(!Xd_0__inst_r_sum1_10__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__9__q ),
	.datab(!Xd_0__inst_r_sum1_8__9__q ),
	.datac(!Xd_0__inst_r_sum1_9__10__q ),
	.datad(!Xd_0__inst_r_sum1_8__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__9__q ),
	.datab(!Xd_0__inst_r_sum1_6__9__q ),
	.datac(!Xd_0__inst_r_sum1_7__10__q ),
	.datad(!Xd_0__inst_r_sum1_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__9__q ),
	.datab(!Xd_0__inst_r_sum1_4__9__q ),
	.datac(!Xd_0__inst_r_sum1_5__10__q ),
	.datad(!Xd_0__inst_r_sum1_4__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__9__q ),
	.datab(!Xd_0__inst_r_sum1_2__9__q ),
	.datac(!Xd_0__inst_r_sum1_3__10__q ),
	.datad(!Xd_0__inst_r_sum1_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__9__q ),
	.datab(!Xd_0__inst_r_sum1_0__9__q ),
	.datac(!Xd_0__inst_r_sum1_1__10__q ),
	.datad(!Xd_0__inst_r_sum1_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__11__q ),
	.datab(!Xd_0__inst_r_sum1_14__11__q ),
	.datac(!Xd_0__inst_r_sum1_14__10__q ),
	.datad(!Xd_0__inst_r_sum1_15__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__11__q ),
	.datab(!Xd_0__inst_r_sum1_12__11__q ),
	.datac(!Xd_0__inst_r_sum1_12__10__q ),
	.datad(!Xd_0__inst_r_sum1_13__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__11__q ),
	.datab(!Xd_0__inst_r_sum1_10__11__q ),
	.datac(!Xd_0__inst_r_sum1_10__10__q ),
	.datad(!Xd_0__inst_r_sum1_11__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__11__q ),
	.datab(!Xd_0__inst_r_sum1_8__11__q ),
	.datac(!Xd_0__inst_r_sum1_8__10__q ),
	.datad(!Xd_0__inst_r_sum1_9__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__11__q ),
	.datab(!Xd_0__inst_r_sum1_6__11__q ),
	.datac(!Xd_0__inst_r_sum1_6__10__q ),
	.datad(!Xd_0__inst_r_sum1_7__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__11__q ),
	.datab(!Xd_0__inst_r_sum1_4__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__10__q ),
	.datad(!Xd_0__inst_r_sum1_5__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__11__q ),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_2__10__q ),
	.datad(!Xd_0__inst_r_sum1_3__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__11__q ),
	.datab(!Xd_0__inst_r_sum1_0__11__q ),
	.datac(!Xd_0__inst_r_sum1_0__10__q ),
	.datad(!Xd_0__inst_r_sum1_1__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__11__q ),
	.datab(!Xd_0__inst_r_sum1_14__11__q ),
	.datac(!Xd_0__inst_r_sum1_15__12__q ),
	.datad(!Xd_0__inst_r_sum1_14__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__11__q ),
	.datab(!Xd_0__inst_r_sum1_12__11__q ),
	.datac(!Xd_0__inst_r_sum1_13__12__q ),
	.datad(!Xd_0__inst_r_sum1_12__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__11__q ),
	.datab(!Xd_0__inst_r_sum1_10__11__q ),
	.datac(!Xd_0__inst_r_sum1_11__12__q ),
	.datad(!Xd_0__inst_r_sum1_10__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__11__q ),
	.datab(!Xd_0__inst_r_sum1_8__11__q ),
	.datac(!Xd_0__inst_r_sum1_9__12__q ),
	.datad(!Xd_0__inst_r_sum1_8__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__11__q ),
	.datab(!Xd_0__inst_r_sum1_6__11__q ),
	.datac(!Xd_0__inst_r_sum1_7__12__q ),
	.datad(!Xd_0__inst_r_sum1_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__11__q ),
	.datab(!Xd_0__inst_r_sum1_4__11__q ),
	.datac(!Xd_0__inst_r_sum1_5__12__q ),
	.datad(!Xd_0__inst_r_sum1_4__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__11__q ),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_3__12__q ),
	.datad(!Xd_0__inst_r_sum1_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__11__q ),
	.datab(!Xd_0__inst_r_sum1_0__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__12__q ),
	.datad(!Xd_0__inst_r_sum1_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__13__q ),
	.datab(!Xd_0__inst_r_sum1_14__13__q ),
	.datac(!Xd_0__inst_r_sum1_14__12__q ),
	.datad(!Xd_0__inst_r_sum1_15__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__13__q ),
	.datab(!Xd_0__inst_r_sum1_12__13__q ),
	.datac(!Xd_0__inst_r_sum1_12__12__q ),
	.datad(!Xd_0__inst_r_sum1_13__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__13__q ),
	.datab(!Xd_0__inst_r_sum1_10__13__q ),
	.datac(!Xd_0__inst_r_sum1_10__12__q ),
	.datad(!Xd_0__inst_r_sum1_11__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__13__q ),
	.datab(!Xd_0__inst_r_sum1_8__13__q ),
	.datac(!Xd_0__inst_r_sum1_8__12__q ),
	.datad(!Xd_0__inst_r_sum1_9__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__13__q ),
	.datab(!Xd_0__inst_r_sum1_6__13__q ),
	.datac(!Xd_0__inst_r_sum1_6__12__q ),
	.datad(!Xd_0__inst_r_sum1_7__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__13__q ),
	.datab(!Xd_0__inst_r_sum1_4__13__q ),
	.datac(!Xd_0__inst_r_sum1_4__12__q ),
	.datad(!Xd_0__inst_r_sum1_5__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__13__q ),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_2__12__q ),
	.datad(!Xd_0__inst_r_sum1_3__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__13__q ),
	.datab(!Xd_0__inst_r_sum1_0__13__q ),
	.datac(!Xd_0__inst_r_sum1_0__12__q ),
	.datad(!Xd_0__inst_r_sum1_1__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__13__q ),
	.datab(!Xd_0__inst_r_sum1_14__13__q ),
	.datac(!Xd_0__inst_r_sum1_15__14__q ),
	.datad(!Xd_0__inst_r_sum1_14__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__13__q ),
	.datab(!Xd_0__inst_r_sum1_12__13__q ),
	.datac(!Xd_0__inst_r_sum1_13__14__q ),
	.datad(!Xd_0__inst_r_sum1_12__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__13__q ),
	.datab(!Xd_0__inst_r_sum1_10__13__q ),
	.datac(!Xd_0__inst_r_sum1_11__14__q ),
	.datad(!Xd_0__inst_r_sum1_10__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__13__q ),
	.datab(!Xd_0__inst_r_sum1_8__13__q ),
	.datac(!Xd_0__inst_r_sum1_9__14__q ),
	.datad(!Xd_0__inst_r_sum1_8__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__13__q ),
	.datab(!Xd_0__inst_r_sum1_6__13__q ),
	.datac(!Xd_0__inst_r_sum1_7__14__q ),
	.datad(!Xd_0__inst_r_sum1_6__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__13__q ),
	.datab(!Xd_0__inst_r_sum1_4__13__q ),
	.datac(!Xd_0__inst_r_sum1_5__14__q ),
	.datad(!Xd_0__inst_r_sum1_4__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__13__q ),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_3__14__q ),
	.datad(!Xd_0__inst_r_sum1_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__13__q ),
	.datab(!Xd_0__inst_r_sum1_0__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__14__q ),
	.datad(!Xd_0__inst_r_sum1_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__15__q ),
	.datab(!Xd_0__inst_r_sum1_15__15__q ),
	.datac(!Xd_0__inst_r_sum1_14__14__q ),
	.datad(!Xd_0__inst_r_sum1_15__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__15__q ),
	.datab(!Xd_0__inst_r_sum1_13__15__q ),
	.datac(!Xd_0__inst_r_sum1_12__14__q ),
	.datad(!Xd_0__inst_r_sum1_13__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__15__q ),
	.datab(!Xd_0__inst_r_sum1_11__15__q ),
	.datac(!Xd_0__inst_r_sum1_10__14__q ),
	.datad(!Xd_0__inst_r_sum1_11__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__15__q ),
	.datab(!Xd_0__inst_r_sum1_9__15__q ),
	.datac(!Xd_0__inst_r_sum1_8__14__q ),
	.datad(!Xd_0__inst_r_sum1_9__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__15__q ),
	.datab(!Xd_0__inst_r_sum1_7__15__q ),
	.datac(!Xd_0__inst_r_sum1_6__14__q ),
	.datad(!Xd_0__inst_r_sum1_7__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__15__q ),
	.datab(!Xd_0__inst_r_sum1_5__15__q ),
	.datac(!Xd_0__inst_r_sum1_4__14__q ),
	.datad(!Xd_0__inst_r_sum1_5__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__15__q ),
	.datab(!Xd_0__inst_r_sum1_3__15__q ),
	.datac(!Xd_0__inst_r_sum1_2__14__q ),
	.datad(!Xd_0__inst_r_sum1_3__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__15__q ),
	.datab(!Xd_0__inst_r_sum1_1__15__q ),
	.datac(!Xd_0__inst_r_sum1_0__14__q ),
	.datad(!Xd_0__inst_r_sum1_1__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__15__q ),
	.datab(!Xd_0__inst_r_sum1_15__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__15__q ),
	.datab(!Xd_0__inst_r_sum1_13__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__15__q ),
	.datab(!Xd_0__inst_r_sum1_11__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__15__q ),
	.datab(!Xd_0__inst_r_sum1_9__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__15__q ),
	.datab(!Xd_0__inst_r_sum1_7__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__15__q ),
	.datab(!Xd_0__inst_r_sum1_5__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__15__q ),
	.datab(!Xd_0__inst_r_sum1_3__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__15__q ),
	.datab(!Xd_0__inst_r_sum1_1__15__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_81_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [12]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [8]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [0]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_87_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [30]),
	.datab(!Xd_0__inst_sign [31]),
	.datac(!Xd_0__inst_product_31__0__q ),
	.datad(!Xd_0__inst_product_30__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [28]),
	.datab(!Xd_0__inst_sign [29]),
	.datac(!Xd_0__inst_product_29__0__q ),
	.datad(!Xd_0__inst_product_28__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_23 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[229]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_23_sumout ),
	.cout(Xd_0__inst_mult_28_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [26]),
	.datab(!Xd_0__inst_sign [27]),
	.datac(!Xd_0__inst_product_27__0__q ),
	.datad(!Xd_0__inst_product_26__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [24]),
	.datab(!Xd_0__inst_sign [25]),
	.datac(!Xd_0__inst_product_25__0__q ),
	.datad(!Xd_0__inst_product_24__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_23 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[245]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_23_sumout ),
	.cout(Xd_0__inst_mult_30_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [22]),
	.datab(!Xd_0__inst_sign [23]),
	.datac(!Xd_0__inst_product_23__0__q ),
	.datad(!Xd_0__inst_product_22__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [20]),
	.datab(!Xd_0__inst_sign [21]),
	.datac(!Xd_0__inst_product_21__0__q ),
	.datad(!Xd_0__inst_product_20__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_23 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[189]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_23_sumout ),
	.cout(Xd_0__inst_mult_23_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [18]),
	.datab(!Xd_0__inst_sign [19]),
	.datac(!Xd_0__inst_product_19__0__q ),
	.datad(!Xd_0__inst_product_18__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [16]),
	.datab(!Xd_0__inst_sign [17]),
	.datac(!Xd_0__inst_product_17__0__q ),
	.datad(!Xd_0__inst_product_16__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_23 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[21]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_23_sumout ),
	.cout(Xd_0__inst_mult_2_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [14]),
	.datab(!Xd_0__inst_sign [15]),
	.datac(!Xd_0__inst_product_15__0__q ),
	.datad(!Xd_0__inst_product_14__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [12]),
	.datab(!Xd_0__inst_sign [13]),
	.datac(!Xd_0__inst_product_13__0__q ),
	.datad(!Xd_0__inst_product_12__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_23 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[37]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_23_sumout ),
	.cout(Xd_0__inst_mult_4_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [10]),
	.datab(!Xd_0__inst_sign [11]),
	.datac(!Xd_0__inst_product_11__0__q ),
	.datad(!Xd_0__inst_product_10__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [8]),
	.datab(!Xd_0__inst_sign [9]),
	.datac(!Xd_0__inst_product_9__0__q ),
	.datad(!Xd_0__inst_product_8__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_23 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[53]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_23_sumout ),
	.cout(Xd_0__inst_mult_6_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [6]),
	.datab(!Xd_0__inst_sign [7]),
	.datac(!Xd_0__inst_product_7__0__q ),
	.datad(!Xd_0__inst_product_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [4]),
	.datab(!Xd_0__inst_sign [5]),
	.datac(!Xd_0__inst_product_5__0__q ),
	.datad(!Xd_0__inst_product_4__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_23 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_23_sumout ),
	.cout(Xd_0__inst_mult_8_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [2]),
	.datab(!Xd_0__inst_sign [3]),
	.datac(!Xd_0__inst_product_3__0__q ),
	.datad(!Xd_0__inst_product_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [0]),
	.datab(!Xd_0__inst_sign [1]),
	.datac(!Xd_0__inst_product_1__0__q ),
	.datad(!Xd_0__inst_product_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_23 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[77]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_23_sumout ),
	.cout(Xd_0__inst_mult_9_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__1__q ),
	.datad(!Xd_0__inst_product_30__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__1__q ),
	.datad(!Xd_0__inst_product_28__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__1__q ),
	.datad(!Xd_0__inst_product_26__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__1__q ),
	.datad(!Xd_0__inst_product_24__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__1__q ),
	.datad(!Xd_0__inst_product_22__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__1__q ),
	.datad(!Xd_0__inst_product_20__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__1__q ),
	.datad(!Xd_0__inst_product_18__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__1__q ),
	.datad(!Xd_0__inst_product_16__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__1__q ),
	.datad(!Xd_0__inst_product_14__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__1__q ),
	.datad(!Xd_0__inst_product_12__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__1__q ),
	.datad(!Xd_0__inst_product_10__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__1__q ),
	.datad(!Xd_0__inst_product_8__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__1__q ),
	.datad(!Xd_0__inst_product_6__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__1__q ),
	.datad(!Xd_0__inst_product_4__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__1__q ),
	.datad(!Xd_0__inst_product_2__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__1__q ),
	.datad(!Xd_0__inst_product_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__2__q ),
	.datad(!Xd_0__inst_product_30__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__2__q ),
	.datad(!Xd_0__inst_product_28__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__2__q ),
	.datad(!Xd_0__inst_product_26__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__2__q ),
	.datad(!Xd_0__inst_product_24__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__2__q ),
	.datad(!Xd_0__inst_product_22__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__2__q ),
	.datad(!Xd_0__inst_product_20__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__2__q ),
	.datad(!Xd_0__inst_product_18__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__2__q ),
	.datad(!Xd_0__inst_product_16__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__2__q ),
	.datad(!Xd_0__inst_product_14__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__2__q ),
	.datad(!Xd_0__inst_product_12__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__2__q ),
	.datad(!Xd_0__inst_product_10__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__2__q ),
	.datad(!Xd_0__inst_product_8__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__2__q ),
	.datad(!Xd_0__inst_product_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__2__q ),
	.datad(!Xd_0__inst_product_4__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__2__q ),
	.datad(!Xd_0__inst_product_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__2__q ),
	.datad(!Xd_0__inst_product_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__3__q ),
	.datad(!Xd_0__inst_product_30__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__3__q ),
	.datad(!Xd_0__inst_product_28__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__3__q ),
	.datad(!Xd_0__inst_product_26__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__3__q ),
	.datad(!Xd_0__inst_product_24__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__3__q ),
	.datad(!Xd_0__inst_product_22__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__3__q ),
	.datad(!Xd_0__inst_product_20__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__3__q ),
	.datad(!Xd_0__inst_product_18__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__3__q ),
	.datad(!Xd_0__inst_product_16__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__3__q ),
	.datad(!Xd_0__inst_product_14__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__3__q ),
	.datad(!Xd_0__inst_product_12__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__3__q ),
	.datad(!Xd_0__inst_product_10__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__3__q ),
	.datad(!Xd_0__inst_product_8__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__3__q ),
	.datad(!Xd_0__inst_product_6__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__3__q ),
	.datad(!Xd_0__inst_product_4__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__3__q ),
	.datad(!Xd_0__inst_product_2__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__3__q ),
	.datad(!Xd_0__inst_product_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__4__q ),
	.datad(!Xd_0__inst_product_30__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__4__q ),
	.datad(!Xd_0__inst_product_28__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__4__q ),
	.datad(!Xd_0__inst_product_26__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__4__q ),
	.datad(!Xd_0__inst_product_24__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__4__q ),
	.datad(!Xd_0__inst_product_22__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__4__q ),
	.datad(!Xd_0__inst_product_20__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__4__q ),
	.datad(!Xd_0__inst_product_18__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__4__q ),
	.datad(!Xd_0__inst_product_16__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__4__q ),
	.datad(!Xd_0__inst_product_14__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__4__q ),
	.datad(!Xd_0__inst_product_12__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__4__q ),
	.datad(!Xd_0__inst_product_10__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__4__q ),
	.datad(!Xd_0__inst_product_8__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__4__q ),
	.datad(!Xd_0__inst_product_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__4__q ),
	.datad(!Xd_0__inst_product_4__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__4__q ),
	.datad(!Xd_0__inst_product_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__4__q ),
	.datad(!Xd_0__inst_product_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__5__q ),
	.datad(!Xd_0__inst_product_30__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__5__q ),
	.datad(!Xd_0__inst_product_28__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__5__q ),
	.datad(!Xd_0__inst_product_26__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__5__q ),
	.datad(!Xd_0__inst_product_24__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__5__q ),
	.datad(!Xd_0__inst_product_22__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__5__q ),
	.datad(!Xd_0__inst_product_20__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__5__q ),
	.datad(!Xd_0__inst_product_18__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__5__q ),
	.datad(!Xd_0__inst_product_16__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__5__q ),
	.datad(!Xd_0__inst_product_14__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__5__q ),
	.datad(!Xd_0__inst_product_12__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__5__q ),
	.datad(!Xd_0__inst_product_10__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__5__q ),
	.datad(!Xd_0__inst_product_8__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__5__q ),
	.datad(!Xd_0__inst_product_6__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__5__q ),
	.datad(!Xd_0__inst_product_4__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__5__q ),
	.datad(!Xd_0__inst_product_2__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__5__q ),
	.datad(!Xd_0__inst_product_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__6__q ),
	.datad(!Xd_0__inst_product_30__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__6__q ),
	.datad(!Xd_0__inst_product_28__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__6__q ),
	.datad(!Xd_0__inst_product_26__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__6__q ),
	.datad(!Xd_0__inst_product_24__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__6__q ),
	.datad(!Xd_0__inst_product_22__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__6__q ),
	.datad(!Xd_0__inst_product_20__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__6__q ),
	.datad(!Xd_0__inst_product_18__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__6__q ),
	.datad(!Xd_0__inst_product_16__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__6__q ),
	.datad(!Xd_0__inst_product_14__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__6__q ),
	.datad(!Xd_0__inst_product_12__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__6__q ),
	.datad(!Xd_0__inst_product_10__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__6__q ),
	.datad(!Xd_0__inst_product_8__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__6__q ),
	.datad(!Xd_0__inst_product_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__6__q ),
	.datad(!Xd_0__inst_product_4__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__6__q ),
	.datad(!Xd_0__inst_product_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__6__q ),
	.datad(!Xd_0__inst_product_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__7__q ),
	.datad(!Xd_0__inst_product_30__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__7__q ),
	.datad(!Xd_0__inst_product_28__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__7__q ),
	.datad(!Xd_0__inst_product_26__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__7__q ),
	.datad(!Xd_0__inst_product_24__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__7__q ),
	.datad(!Xd_0__inst_product_22__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__7__q ),
	.datad(!Xd_0__inst_product_20__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__7__q ),
	.datad(!Xd_0__inst_product_18__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__7__q ),
	.datad(!Xd_0__inst_product_16__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__7__q ),
	.datad(!Xd_0__inst_product_14__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__7__q ),
	.datad(!Xd_0__inst_product_12__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__7__q ),
	.datad(!Xd_0__inst_product_10__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__7__q ),
	.datad(!Xd_0__inst_product_8__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__7__q ),
	.datad(!Xd_0__inst_product_6__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__7__q ),
	.datad(!Xd_0__inst_product_4__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__7__q ),
	.datad(!Xd_0__inst_product_2__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__7__q ),
	.datad(!Xd_0__inst_product_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__8__q ),
	.datad(!Xd_0__inst_product_30__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__8__q ),
	.datad(!Xd_0__inst_product_28__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__8__q ),
	.datad(!Xd_0__inst_product_26__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__8__q ),
	.datad(!Xd_0__inst_product_24__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__8__q ),
	.datad(!Xd_0__inst_product_22__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__8__q ),
	.datad(!Xd_0__inst_product_20__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__8__q ),
	.datad(!Xd_0__inst_product_18__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__8__q ),
	.datad(!Xd_0__inst_product_16__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__8__q ),
	.datad(!Xd_0__inst_product_14__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__8__q ),
	.datad(!Xd_0__inst_product_12__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__8__q ),
	.datad(!Xd_0__inst_product_10__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__8__q ),
	.datad(!Xd_0__inst_product_8__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__8__q ),
	.datad(!Xd_0__inst_product_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__8__q ),
	.datad(!Xd_0__inst_product_4__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__8__q ),
	.datad(!Xd_0__inst_product_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__8__q ),
	.datad(!Xd_0__inst_product_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__9__q ),
	.datad(!Xd_0__inst_product_30__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__9__q ),
	.datad(!Xd_0__inst_product_28__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__9__q ),
	.datad(!Xd_0__inst_product_26__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__9__q ),
	.datad(!Xd_0__inst_product_24__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__9__q ),
	.datad(!Xd_0__inst_product_22__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__9__q ),
	.datad(!Xd_0__inst_product_20__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__9__q ),
	.datad(!Xd_0__inst_product_18__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__9__q ),
	.datad(!Xd_0__inst_product_16__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__9__q ),
	.datad(!Xd_0__inst_product_14__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__9__q ),
	.datad(!Xd_0__inst_product_12__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__9__q ),
	.datad(!Xd_0__inst_product_10__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__9__q ),
	.datad(!Xd_0__inst_product_8__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__9__q ),
	.datad(!Xd_0__inst_product_6__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__9__q ),
	.datad(!Xd_0__inst_product_4__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__9__q ),
	.datad(!Xd_0__inst_product_2__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__9__q ),
	.datad(!Xd_0__inst_product_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__10__q ),
	.datad(!Xd_0__inst_product_30__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__10__q ),
	.datad(!Xd_0__inst_product_28__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__10__q ),
	.datad(!Xd_0__inst_product_26__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__10__q ),
	.datad(!Xd_0__inst_product_24__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__10__q ),
	.datad(!Xd_0__inst_product_22__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__10__q ),
	.datad(!Xd_0__inst_product_20__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__10__q ),
	.datad(!Xd_0__inst_product_18__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__10__q ),
	.datad(!Xd_0__inst_product_16__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__10__q ),
	.datad(!Xd_0__inst_product_14__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__10__q ),
	.datad(!Xd_0__inst_product_12__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__10__q ),
	.datad(!Xd_0__inst_product_10__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__10__q ),
	.datad(!Xd_0__inst_product_8__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__10__q ),
	.datad(!Xd_0__inst_product_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__10__q ),
	.datad(!Xd_0__inst_product_4__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__10__q ),
	.datad(!Xd_0__inst_product_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__10__q ),
	.datad(!Xd_0__inst_product_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__11__q ),
	.datad(!Xd_0__inst_product_30__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__11__q ),
	.datad(!Xd_0__inst_product_28__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__11__q ),
	.datad(!Xd_0__inst_product_26__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__11__q ),
	.datad(!Xd_0__inst_product_24__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__11__q ),
	.datad(!Xd_0__inst_product_22__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__11__q ),
	.datad(!Xd_0__inst_product_20__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__11__q ),
	.datad(!Xd_0__inst_product_18__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__11__q ),
	.datad(!Xd_0__inst_product_16__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__11__q ),
	.datad(!Xd_0__inst_product_14__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__11__q ),
	.datad(!Xd_0__inst_product_12__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__11__q ),
	.datad(!Xd_0__inst_product_10__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__11__q ),
	.datad(!Xd_0__inst_product_8__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__11__q ),
	.datad(!Xd_0__inst_product_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__11__q ),
	.datad(!Xd_0__inst_product_4__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__11__q ),
	.datad(!Xd_0__inst_product_2__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__11__q ),
	.datad(!Xd_0__inst_product_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__12__q ),
	.datad(!Xd_0__inst_product_30__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__12__q ),
	.datad(!Xd_0__inst_product_28__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__12__q ),
	.datad(!Xd_0__inst_product_26__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__12__q ),
	.datad(!Xd_0__inst_product_24__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__12__q ),
	.datad(!Xd_0__inst_product_22__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__12__q ),
	.datad(!Xd_0__inst_product_20__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__12__q ),
	.datad(!Xd_0__inst_product_18__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__12__q ),
	.datad(!Xd_0__inst_product_16__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__12__q ),
	.datad(!Xd_0__inst_product_14__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__12__q ),
	.datad(!Xd_0__inst_product_12__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__12__q ),
	.datad(!Xd_0__inst_product_10__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__12__q ),
	.datad(!Xd_0__inst_product_8__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__12__q ),
	.datad(!Xd_0__inst_product_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__12__q ),
	.datad(!Xd_0__inst_product_4__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__12__q ),
	.datad(!Xd_0__inst_product_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__12__q ),
	.datad(!Xd_0__inst_product_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__13__q ),
	.datad(!Xd_0__inst_product_30__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__13__q ),
	.datad(!Xd_0__inst_product_28__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__13__q ),
	.datad(!Xd_0__inst_product_26__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__13__q ),
	.datad(!Xd_0__inst_product_24__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__13__q ),
	.datad(!Xd_0__inst_product_22__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__13__q ),
	.datad(!Xd_0__inst_product_20__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__13__q ),
	.datad(!Xd_0__inst_product_18__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__13__q ),
	.datad(!Xd_0__inst_product_16__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__13__q ),
	.datad(!Xd_0__inst_product_14__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__13__q ),
	.datad(!Xd_0__inst_product_12__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__13__q ),
	.datad(!Xd_0__inst_product_10__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__13__q ),
	.datad(!Xd_0__inst_product_8__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__13__q ),
	.datad(!Xd_0__inst_product_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__13__q ),
	.datad(!Xd_0__inst_product_4__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__13__q ),
	.datad(!Xd_0__inst_product_2__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__13__q ),
	.datad(!Xd_0__inst_product_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [29]),
	.datad(!Xd_0__inst_sign [28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [31]),
	.datad(!Xd_0__inst_sign [30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [25]),
	.datad(!Xd_0__inst_sign [24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [27]),
	.datad(!Xd_0__inst_sign [26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [21]),
	.datad(!Xd_0__inst_sign [20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [23]),
	.datad(!Xd_0__inst_sign [22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [17]),
	.datad(!Xd_0__inst_sign [16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [19]),
	.datad(!Xd_0__inst_sign [18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [13]),
	.datad(!Xd_0__inst_sign [12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [15]),
	.datad(!Xd_0__inst_sign [14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [9]),
	.datad(!Xd_0__inst_sign [8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [11]),
	.datad(!Xd_0__inst_sign [10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [5]),
	.datad(!Xd_0__inst_sign [4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [7]),
	.datad(!Xd_0__inst_sign [6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [1]),
	.datad(!Xd_0__inst_sign [0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [3]),
	.datad(!Xd_0__inst_sign [2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_76_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [30]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [28]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_23 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[221]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_23_sumout ),
	.cout(Xd_0__inst_mult_27_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [26]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [24]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_23 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[237]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_23_sumout ),
	.cout(Xd_0__inst_mult_29_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [22]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [20]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_28 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[86]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_28_sumout ),
	.cout(Xd_0__inst_mult_10_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [18]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [16]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_23 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[253]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_23_sumout ),
	.cout(Xd_0__inst_mult_31_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [14]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [12]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_23 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[29]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_23_sumout ),
	.cout(Xd_0__inst_mult_3_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [10]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [8]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_23 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[45]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_23_sumout ),
	.cout(Xd_0__inst_mult_5_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [6]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_23 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[61]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_23_sumout ),
	.cout(Xd_0__inst_mult_7_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_85 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_23 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[13]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_23_sumout ),
	.cout(Xd_0__inst_mult_1_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_83 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[43]),
	.datac(!din_a[44]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_84 ),
	.cout(Xd_0__inst_mult_5_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_83 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[51]),
	.datac(!din_a[52]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_84 ),
	.cout(Xd_0__inst_mult_6_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_1 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[255]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_1_sumout ),
	.cout(Xd_0__inst_i21_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_83 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[59]),
	.datac(!din_a[60]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_84 ),
	.cout(Xd_0__inst_mult_7_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_83 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[67]),
	.datac(!din_a[68]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_84 ),
	.cout(Xd_0__inst_mult_8_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_6 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[223]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_6_sumout ),
	.cout(Xd_0__inst_i21_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_83 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[75]),
	.datac(!din_a[76]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_84 ),
	.cout(Xd_0__inst_mult_9_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_83 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[163]),
	.datac(!din_a[164]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_84 ),
	.cout(Xd_0__inst_mult_20_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_11 (
// Equation(s):

	.dataa(!din_a[191]),
	.datab(!din_b[191]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_11_sumout ),
	.cout(Xd_0__inst_i21_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_83 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[155]),
	.datac(!din_a[156]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_84 ),
	.cout(Xd_0__inst_mult_19_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_83 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[91]),
	.datac(!din_a[92]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_84 ),
	.cout(Xd_0__inst_mult_11_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_16 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[159]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_16_sumout ),
	.cout(Xd_0__inst_i21_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_83 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[147]),
	.datac(!din_a[148]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_84 ),
	.cout(Xd_0__inst_mult_18_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_83 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[139]),
	.datac(!din_a[140]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_84 ),
	.cout(Xd_0__inst_mult_17_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_21 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[127]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_21_sumout ),
	.cout(Xd_0__inst_i21_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_83 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[131]),
	.datac(!din_a[132]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_84 ),
	.cout(Xd_0__inst_mult_16_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_83 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[83]),
	.datac(!din_a[84]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_84 ),
	.cout(Xd_0__inst_mult_10_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_26 (
// Equation(s):

	.dataa(!din_a[95]),
	.datab(!din_b[95]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_26_sumout ),
	.cout(Xd_0__inst_i21_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_83 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[123]),
	.datac(!din_a[124]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_84 ),
	.cout(Xd_0__inst_mult_15_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_83 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[115]),
	.datac(!din_a[116]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_84 ),
	.cout(Xd_0__inst_mult_14_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_31 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[63]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_31_sumout ),
	.cout(Xd_0__inst_i21_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_83 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[107]),
	.datac(!din_a[108]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_84 ),
	.cout(Xd_0__inst_mult_13_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_83 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[99]),
	.datac(!din_a[100]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_84 ),
	.cout(Xd_0__inst_mult_12_85 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_36 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_36_sumout ),
	.cout(Xd_0__inst_i21_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_0_q ),
	.datab(!Xd_0__inst_mult_31_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_85 ),
	.cout(Xd_0__inst_mult_31_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_0_q ),
	.datab(!Xd_0__inst_mult_30_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_85 ),
	.cout(Xd_0__inst_mult_30_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_0_q ),
	.datab(!Xd_0__inst_mult_29_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_85 ),
	.cout(Xd_0__inst_mult_29_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_0_q ),
	.datab(!Xd_0__inst_mult_28_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_85 ),
	.cout(Xd_0__inst_mult_28_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_0_q ),
	.datab(!Xd_0__inst_mult_27_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_85 ),
	.cout(Xd_0__inst_mult_27_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_0_q ),
	.datab(!Xd_0__inst_mult_26_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_85 ),
	.cout(Xd_0__inst_mult_26_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_0_q ),
	.datab(!Xd_0__inst_mult_25_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_85 ),
	.cout(Xd_0__inst_mult_25_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_0_q ),
	.datab(!Xd_0__inst_mult_24_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_85 ),
	.cout(Xd_0__inst_mult_24_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_0_q ),
	.datab(!Xd_0__inst_mult_23_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_85 ),
	.cout(Xd_0__inst_mult_23_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_0_q ),
	.datab(!Xd_0__inst_mult_22_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_85 ),
	.cout(Xd_0__inst_mult_22_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_0_q ),
	.datab(!Xd_0__inst_mult_21_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_85 ),
	.cout(Xd_0__inst_mult_21_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_0_q ),
	.datab(!Xd_0__inst_mult_20_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_89 ),
	.cout(Xd_0__inst_mult_20_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_0_q ),
	.datab(!Xd_0__inst_mult_19_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_89 ),
	.cout(Xd_0__inst_mult_19_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_0_q ),
	.datab(!Xd_0__inst_mult_18_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_89 ),
	.cout(Xd_0__inst_mult_18_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_0_q ),
	.datab(!Xd_0__inst_mult_17_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_89 ),
	.cout(Xd_0__inst_mult_17_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_0_q ),
	.datab(!Xd_0__inst_mult_16_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_89 ),
	.cout(Xd_0__inst_mult_16_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_0_q ),
	.datab(!Xd_0__inst_mult_15_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_89 ),
	.cout(Xd_0__inst_mult_15_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_0_q ),
	.datab(!Xd_0__inst_mult_14_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_89 ),
	.cout(Xd_0__inst_mult_14_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_0_q ),
	.datab(!Xd_0__inst_mult_13_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_89 ),
	.cout(Xd_0__inst_mult_13_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_0_q ),
	.datab(!Xd_0__inst_mult_12_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_89 ),
	.cout(Xd_0__inst_mult_12_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_0_q ),
	.datab(!Xd_0__inst_mult_11_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_89 ),
	.cout(Xd_0__inst_mult_11_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_0_q ),
	.datab(!Xd_0__inst_mult_10_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_89 ),
	.cout(Xd_0__inst_mult_10_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_0_q ),
	.datab(!Xd_0__inst_mult_9_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_89 ),
	.cout(Xd_0__inst_mult_9_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_0_q ),
	.datab(!Xd_0__inst_mult_8_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_89 ),
	.cout(Xd_0__inst_mult_8_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_164 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_89 ),
	.cout(Xd_0__inst_mult_7_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_89 ),
	.cout(Xd_0__inst_mult_6_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_89 ),
	.cout(Xd_0__inst_mult_5_90 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_85 ),
	.cout(Xd_0__inst_mult_4_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_0_q ),
	.datab(!Xd_0__inst_mult_3_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_85 ),
	.cout(Xd_0__inst_mult_3_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_0_q ),
	.datab(!Xd_0__inst_mult_2_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_85 ),
	.cout(Xd_0__inst_mult_2_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_0_q ),
	.datab(!Xd_0__inst_mult_1_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_85 ),
	.cout(Xd_0__inst_mult_1_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_0_q ),
	.datab(!Xd_0__inst_mult_0_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_85 ),
	.cout(Xd_0__inst_mult_0_86 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_2_q ),
	.datab(!Xd_0__inst_mult_31_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_90 ),
	.cout(Xd_0__inst_mult_31_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_2_q ),
	.datab(!Xd_0__inst_mult_30_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_90 ),
	.cout(Xd_0__inst_mult_30_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_2_q ),
	.datab(!Xd_0__inst_mult_29_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_90 ),
	.cout(Xd_0__inst_mult_29_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_2_q ),
	.datab(!Xd_0__inst_mult_28_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_90 ),
	.cout(Xd_0__inst_mult_28_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_2_q ),
	.datab(!Xd_0__inst_mult_27_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_90 ),
	.cout(Xd_0__inst_mult_27_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_2_q ),
	.datab(!Xd_0__inst_mult_26_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_90 ),
	.cout(Xd_0__inst_mult_26_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_2_q ),
	.datab(!Xd_0__inst_mult_25_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_90 ),
	.cout(Xd_0__inst_mult_25_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_2_q ),
	.datab(!Xd_0__inst_mult_24_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_90 ),
	.cout(Xd_0__inst_mult_24_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_2_q ),
	.datab(!Xd_0__inst_mult_23_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_90 ),
	.cout(Xd_0__inst_mult_23_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_2_q ),
	.datab(!Xd_0__inst_mult_22_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_90 ),
	.cout(Xd_0__inst_mult_22_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_2_q ),
	.datab(!Xd_0__inst_mult_21_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_90 ),
	.cout(Xd_0__inst_mult_21_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_2_q ),
	.datab(!Xd_0__inst_mult_20_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_93 ),
	.cout(Xd_0__inst_mult_20_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_2_q ),
	.datab(!Xd_0__inst_mult_19_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_93 ),
	.cout(Xd_0__inst_mult_19_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_2_q ),
	.datab(!Xd_0__inst_mult_18_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_93 ),
	.cout(Xd_0__inst_mult_18_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_2_q ),
	.datab(!Xd_0__inst_mult_17_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_93 ),
	.cout(Xd_0__inst_mult_17_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_2_q ),
	.datab(!Xd_0__inst_mult_16_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_93 ),
	.cout(Xd_0__inst_mult_16_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_2_q ),
	.datab(!Xd_0__inst_mult_15_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_93 ),
	.cout(Xd_0__inst_mult_15_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_2_q ),
	.datab(!Xd_0__inst_mult_14_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_93 ),
	.cout(Xd_0__inst_mult_14_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_2_q ),
	.datab(!Xd_0__inst_mult_13_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_93 ),
	.cout(Xd_0__inst_mult_13_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_2_q ),
	.datab(!Xd_0__inst_mult_12_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_93 ),
	.cout(Xd_0__inst_mult_12_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_2_q ),
	.datab(!Xd_0__inst_mult_11_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_93 ),
	.cout(Xd_0__inst_mult_11_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_2_q ),
	.datab(!Xd_0__inst_mult_10_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_93 ),
	.cout(Xd_0__inst_mult_10_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_2_q ),
	.datab(!Xd_0__inst_mult_9_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_93 ),
	.cout(Xd_0__inst_mult_9_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_2_q ),
	.datab(!Xd_0__inst_mult_8_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_93 ),
	.cout(Xd_0__inst_mult_8_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_2_q ),
	.datab(!Xd_0__inst_mult_7_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_93 ),
	.cout(Xd_0__inst_mult_7_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_2_q ),
	.datab(!Xd_0__inst_mult_6_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_93 ),
	.cout(Xd_0__inst_mult_6_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_2_q ),
	.datab(!Xd_0__inst_mult_5_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_90 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_93 ),
	.cout(Xd_0__inst_mult_5_94 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_2_q ),
	.datab(!Xd_0__inst_mult_4_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_90 ),
	.cout(Xd_0__inst_mult_4_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_2_q ),
	.datab(!Xd_0__inst_mult_3_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_90 ),
	.cout(Xd_0__inst_mult_3_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_2_q ),
	.datab(!Xd_0__inst_mult_2_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_90 ),
	.cout(Xd_0__inst_mult_2_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_2_q ),
	.datab(!Xd_0__inst_mult_1_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_90 ),
	.cout(Xd_0__inst_mult_1_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_2_q ),
	.datab(!Xd_0__inst_mult_0_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_86 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_90 ),
	.cout(Xd_0__inst_mult_0_91 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_4_q ),
	.datab(!Xd_0__inst_mult_31_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_94 ),
	.cout(Xd_0__inst_mult_31_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_4_q ),
	.datab(!Xd_0__inst_mult_30_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_94 ),
	.cout(Xd_0__inst_mult_30_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_4_q ),
	.datab(!Xd_0__inst_mult_29_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_94 ),
	.cout(Xd_0__inst_mult_29_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_4_q ),
	.datab(!Xd_0__inst_mult_28_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_94 ),
	.cout(Xd_0__inst_mult_28_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_4_q ),
	.datab(!Xd_0__inst_mult_27_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_94 ),
	.cout(Xd_0__inst_mult_27_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_4_q ),
	.datab(!Xd_0__inst_mult_26_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_94 ),
	.cout(Xd_0__inst_mult_26_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_4_q ),
	.datab(!Xd_0__inst_mult_25_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_94 ),
	.cout(Xd_0__inst_mult_25_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_4_q ),
	.datab(!Xd_0__inst_mult_24_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_94 ),
	.cout(Xd_0__inst_mult_24_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_4_q ),
	.datab(!Xd_0__inst_mult_23_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_94 ),
	.cout(Xd_0__inst_mult_23_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_4_q ),
	.datab(!Xd_0__inst_mult_22_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_94 ),
	.cout(Xd_0__inst_mult_22_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_4_q ),
	.datab(!Xd_0__inst_mult_21_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_94 ),
	.cout(Xd_0__inst_mult_21_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_4_q ),
	.datab(!Xd_0__inst_mult_20_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_98 ),
	.cout(Xd_0__inst_mult_20_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_4_q ),
	.datab(!Xd_0__inst_mult_19_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_98 ),
	.cout(Xd_0__inst_mult_19_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_4_q ),
	.datab(!Xd_0__inst_mult_18_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_98 ),
	.cout(Xd_0__inst_mult_18_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_4_q ),
	.datab(!Xd_0__inst_mult_17_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_98 ),
	.cout(Xd_0__inst_mult_17_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_4_q ),
	.datab(!Xd_0__inst_mult_16_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_98 ),
	.cout(Xd_0__inst_mult_16_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_98 ),
	.cout(Xd_0__inst_mult_15_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_98 ),
	.cout(Xd_0__inst_mult_14_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_98 ),
	.cout(Xd_0__inst_mult_13_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_98 ),
	.cout(Xd_0__inst_mult_12_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_98 ),
	.cout(Xd_0__inst_mult_11_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_98 ),
	.cout(Xd_0__inst_mult_10_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_98 ),
	.cout(Xd_0__inst_mult_9_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_98 ),
	.cout(Xd_0__inst_mult_8_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_98 ),
	.cout(Xd_0__inst_mult_7_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_98 ),
	.cout(Xd_0__inst_mult_6_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_94 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_98 ),
	.cout(Xd_0__inst_mult_5_99 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_94 ),
	.cout(Xd_0__inst_mult_4_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_94 ),
	.cout(Xd_0__inst_mult_3_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_94 ),
	.cout(Xd_0__inst_mult_2_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_94 ),
	.cout(Xd_0__inst_mult_1_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_37 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_91 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_94 ),
	.cout(Xd_0__inst_mult_0_95 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_6_q ),
	.datab(!Xd_0__inst_mult_31_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_99 ),
	.cout(Xd_0__inst_mult_31_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_6_q ),
	.datab(!Xd_0__inst_mult_30_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_99 ),
	.cout(Xd_0__inst_mult_30_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_6_q ),
	.datab(!Xd_0__inst_mult_29_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_99 ),
	.cout(Xd_0__inst_mult_29_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_6_q ),
	.datab(!Xd_0__inst_mult_28_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_99 ),
	.cout(Xd_0__inst_mult_28_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_6_q ),
	.datab(!Xd_0__inst_mult_27_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_99 ),
	.cout(Xd_0__inst_mult_27_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_6_q ),
	.datab(!Xd_0__inst_mult_26_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_99 ),
	.cout(Xd_0__inst_mult_26_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_6_q ),
	.datab(!Xd_0__inst_mult_25_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_99 ),
	.cout(Xd_0__inst_mult_25_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_6_q ),
	.datab(!Xd_0__inst_mult_24_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_99 ),
	.cout(Xd_0__inst_mult_24_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_6_q ),
	.datab(!Xd_0__inst_mult_23_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_99 ),
	.cout(Xd_0__inst_mult_23_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_6_q ),
	.datab(!Xd_0__inst_mult_22_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_99 ),
	.cout(Xd_0__inst_mult_22_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_6_q ),
	.datab(!Xd_0__inst_mult_21_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_99 ),
	.cout(Xd_0__inst_mult_21_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_6_q ),
	.datab(!Xd_0__inst_mult_20_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_103 ),
	.cout(Xd_0__inst_mult_20_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_6_q ),
	.datab(!Xd_0__inst_mult_19_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_103 ),
	.cout(Xd_0__inst_mult_19_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_6_q ),
	.datab(!Xd_0__inst_mult_18_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_103 ),
	.cout(Xd_0__inst_mult_18_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_6_q ),
	.datab(!Xd_0__inst_mult_17_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_103 ),
	.cout(Xd_0__inst_mult_17_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_6_q ),
	.datab(!Xd_0__inst_mult_16_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_103 ),
	.cout(Xd_0__inst_mult_16_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_6_q ),
	.datab(!Xd_0__inst_mult_15_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_103 ),
	.cout(Xd_0__inst_mult_15_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_6_q ),
	.datab(!Xd_0__inst_mult_14_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_103 ),
	.cout(Xd_0__inst_mult_14_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_6_q ),
	.datab(!Xd_0__inst_mult_13_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_103 ),
	.cout(Xd_0__inst_mult_13_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_6_q ),
	.datab(!Xd_0__inst_mult_12_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_103 ),
	.cout(Xd_0__inst_mult_12_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_6_q ),
	.datab(!Xd_0__inst_mult_11_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_103 ),
	.cout(Xd_0__inst_mult_11_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_6_q ),
	.datab(!Xd_0__inst_mult_10_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_103 ),
	.cout(Xd_0__inst_mult_10_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_6_q ),
	.datab(!Xd_0__inst_mult_9_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_103 ),
	.cout(Xd_0__inst_mult_9_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_6_q ),
	.datab(!Xd_0__inst_mult_8_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_103 ),
	.cout(Xd_0__inst_mult_8_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_6_q ),
	.datab(!Xd_0__inst_mult_7_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_103 ),
	.cout(Xd_0__inst_mult_7_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_6_q ),
	.datab(!Xd_0__inst_mult_6_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_103 ),
	.cout(Xd_0__inst_mult_6_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_6_q ),
	.datab(!Xd_0__inst_mult_5_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_99 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_103 ),
	.cout(Xd_0__inst_mult_5_104 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_6_q ),
	.datab(!Xd_0__inst_mult_4_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_99 ),
	.cout(Xd_0__inst_mult_4_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_6_q ),
	.datab(!Xd_0__inst_mult_3_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_99 ),
	.cout(Xd_0__inst_mult_3_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_6_q ),
	.datab(!Xd_0__inst_mult_2_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_99 ),
	.cout(Xd_0__inst_mult_2_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_6_q ),
	.datab(!Xd_0__inst_mult_1_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_99 ),
	.cout(Xd_0__inst_mult_1_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_38 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_6_q ),
	.datab(!Xd_0__inst_mult_0_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_95 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_99 ),
	.cout(Xd_0__inst_mult_0_100 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_8_q ),
	.datab(!Xd_0__inst_mult_31_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_104 ),
	.cout(Xd_0__inst_mult_31_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_8_q ),
	.datab(!Xd_0__inst_mult_30_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_104 ),
	.cout(Xd_0__inst_mult_30_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_8_q ),
	.datab(!Xd_0__inst_mult_29_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_104 ),
	.cout(Xd_0__inst_mult_29_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_8_q ),
	.datab(!Xd_0__inst_mult_28_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_104 ),
	.cout(Xd_0__inst_mult_28_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_8_q ),
	.datab(!Xd_0__inst_mult_27_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_104 ),
	.cout(Xd_0__inst_mult_27_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_8_q ),
	.datab(!Xd_0__inst_mult_26_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_104 ),
	.cout(Xd_0__inst_mult_26_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_8_q ),
	.datab(!Xd_0__inst_mult_25_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_104 ),
	.cout(Xd_0__inst_mult_25_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_8_q ),
	.datab(!Xd_0__inst_mult_24_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_104 ),
	.cout(Xd_0__inst_mult_24_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_8_q ),
	.datab(!Xd_0__inst_mult_23_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_104 ),
	.cout(Xd_0__inst_mult_23_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_8_q ),
	.datab(!Xd_0__inst_mult_22_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_104 ),
	.cout(Xd_0__inst_mult_22_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_8_q ),
	.datab(!Xd_0__inst_mult_21_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_104 ),
	.cout(Xd_0__inst_mult_21_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_8_q ),
	.datab(!Xd_0__inst_mult_20_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_108 ),
	.cout(Xd_0__inst_mult_20_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_8_q ),
	.datab(!Xd_0__inst_mult_19_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_108 ),
	.cout(Xd_0__inst_mult_19_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_8_q ),
	.datab(!Xd_0__inst_mult_18_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_108 ),
	.cout(Xd_0__inst_mult_18_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_8_q ),
	.datab(!Xd_0__inst_mult_17_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_108 ),
	.cout(Xd_0__inst_mult_17_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_8_q ),
	.datab(!Xd_0__inst_mult_16_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_108 ),
	.cout(Xd_0__inst_mult_16_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_8_q ),
	.datab(!Xd_0__inst_mult_15_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_108 ),
	.cout(Xd_0__inst_mult_15_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_8_q ),
	.datab(!Xd_0__inst_mult_14_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_108 ),
	.cout(Xd_0__inst_mult_14_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_8_q ),
	.datab(!Xd_0__inst_mult_13_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_108 ),
	.cout(Xd_0__inst_mult_13_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_8_q ),
	.datab(!Xd_0__inst_mult_12_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_108 ),
	.cout(Xd_0__inst_mult_12_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_8_q ),
	.datab(!Xd_0__inst_mult_11_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_108 ),
	.cout(Xd_0__inst_mult_11_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_8_q ),
	.datab(!Xd_0__inst_mult_10_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_108 ),
	.cout(Xd_0__inst_mult_10_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_8_q ),
	.datab(!Xd_0__inst_mult_9_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_108 ),
	.cout(Xd_0__inst_mult_9_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_8_q ),
	.datab(!Xd_0__inst_mult_8_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_108 ),
	.cout(Xd_0__inst_mult_8_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_8_q ),
	.datab(!Xd_0__inst_mult_7_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_108 ),
	.cout(Xd_0__inst_mult_7_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_8_q ),
	.datab(!Xd_0__inst_mult_6_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_108 ),
	.cout(Xd_0__inst_mult_6_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_8_q ),
	.datab(!Xd_0__inst_mult_5_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_104 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_108 ),
	.cout(Xd_0__inst_mult_5_109 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_8_q ),
	.datab(!Xd_0__inst_mult_4_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_104 ),
	.cout(Xd_0__inst_mult_4_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_8_q ),
	.datab(!Xd_0__inst_mult_3_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_104 ),
	.cout(Xd_0__inst_mult_3_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_8_q ),
	.datab(!Xd_0__inst_mult_2_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_104 ),
	.cout(Xd_0__inst_mult_2_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_8_q ),
	.datab(!Xd_0__inst_mult_1_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_104 ),
	.cout(Xd_0__inst_mult_1_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_39 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_8_q ),
	.datab(!Xd_0__inst_mult_0_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_100 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_104 ),
	.cout(Xd_0__inst_mult_0_105 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_10_q ),
	.datab(!Xd_0__inst_mult_31_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_109 ),
	.cout(Xd_0__inst_mult_31_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_10_q ),
	.datab(!Xd_0__inst_mult_30_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_109 ),
	.cout(Xd_0__inst_mult_30_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_10_q ),
	.datab(!Xd_0__inst_mult_29_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_109 ),
	.cout(Xd_0__inst_mult_29_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_10_q ),
	.datab(!Xd_0__inst_mult_28_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_109 ),
	.cout(Xd_0__inst_mult_28_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_10_q ),
	.datab(!Xd_0__inst_mult_27_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_109 ),
	.cout(Xd_0__inst_mult_27_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_10_q ),
	.datab(!Xd_0__inst_mult_26_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_109 ),
	.cout(Xd_0__inst_mult_26_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_10_q ),
	.datab(!Xd_0__inst_mult_25_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_109 ),
	.cout(Xd_0__inst_mult_25_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_10_q ),
	.datab(!Xd_0__inst_mult_24_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_109 ),
	.cout(Xd_0__inst_mult_24_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_10_q ),
	.datab(!Xd_0__inst_mult_23_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_109 ),
	.cout(Xd_0__inst_mult_23_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_10_q ),
	.datab(!Xd_0__inst_mult_22_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_109 ),
	.cout(Xd_0__inst_mult_22_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_10_q ),
	.datab(!Xd_0__inst_mult_21_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_109 ),
	.cout(Xd_0__inst_mult_21_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_10_q ),
	.datab(!Xd_0__inst_mult_20_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_113 ),
	.cout(Xd_0__inst_mult_20_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_10_q ),
	.datab(!Xd_0__inst_mult_19_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_113 ),
	.cout(Xd_0__inst_mult_19_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_10_q ),
	.datab(!Xd_0__inst_mult_18_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_113 ),
	.cout(Xd_0__inst_mult_18_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_10_q ),
	.datab(!Xd_0__inst_mult_17_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_113 ),
	.cout(Xd_0__inst_mult_17_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_10_q ),
	.datab(!Xd_0__inst_mult_16_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_113 ),
	.cout(Xd_0__inst_mult_16_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_10_q ),
	.datab(!Xd_0__inst_mult_15_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_113 ),
	.cout(Xd_0__inst_mult_15_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_10_q ),
	.datab(!Xd_0__inst_mult_14_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_113 ),
	.cout(Xd_0__inst_mult_14_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_10_q ),
	.datab(!Xd_0__inst_mult_13_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_113 ),
	.cout(Xd_0__inst_mult_13_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_10_q ),
	.datab(!Xd_0__inst_mult_12_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_113 ),
	.cout(Xd_0__inst_mult_12_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_10_q ),
	.datab(!Xd_0__inst_mult_11_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_113 ),
	.cout(Xd_0__inst_mult_11_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_10_q ),
	.datab(!Xd_0__inst_mult_10_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_113 ),
	.cout(Xd_0__inst_mult_10_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_10_q ),
	.datab(!Xd_0__inst_mult_9_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_113 ),
	.cout(Xd_0__inst_mult_9_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_10_q ),
	.datab(!Xd_0__inst_mult_8_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_113 ),
	.cout(Xd_0__inst_mult_8_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_10_q ),
	.datab(!Xd_0__inst_mult_7_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_113 ),
	.cout(Xd_0__inst_mult_7_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_10_q ),
	.datab(!Xd_0__inst_mult_6_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_113 ),
	.cout(Xd_0__inst_mult_6_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_10_q ),
	.datab(!Xd_0__inst_mult_5_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_109 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_113 ),
	.cout(Xd_0__inst_mult_5_114 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_10_q ),
	.datab(!Xd_0__inst_mult_4_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_109 ),
	.cout(Xd_0__inst_mult_4_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_10_q ),
	.datab(!Xd_0__inst_mult_3_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_109 ),
	.cout(Xd_0__inst_mult_3_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_10_q ),
	.datab(!Xd_0__inst_mult_2_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_109 ),
	.cout(Xd_0__inst_mult_2_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_10_q ),
	.datab(!Xd_0__inst_mult_1_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_109 ),
	.cout(Xd_0__inst_mult_1_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_40 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_10_q ),
	.datab(!Xd_0__inst_mult_0_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_105 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_109 ),
	.cout(Xd_0__inst_mult_0_110 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_12_q ),
	.datab(!Xd_0__inst_mult_31_13_q ),
	.datac(!Xd_0__inst_mult_31_14_q ),
	.datad(!Xd_0__inst_mult_31_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_114 ),
	.cout(Xd_0__inst_mult_31_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_12_q ),
	.datab(!Xd_0__inst_mult_30_13_q ),
	.datac(!Xd_0__inst_mult_30_14_q ),
	.datad(!Xd_0__inst_mult_30_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_114 ),
	.cout(Xd_0__inst_mult_30_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_12_q ),
	.datab(!Xd_0__inst_mult_29_13_q ),
	.datac(!Xd_0__inst_mult_29_14_q ),
	.datad(!Xd_0__inst_mult_29_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_114 ),
	.cout(Xd_0__inst_mult_29_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_12_q ),
	.datab(!Xd_0__inst_mult_28_13_q ),
	.datac(!Xd_0__inst_mult_28_14_q ),
	.datad(!Xd_0__inst_mult_28_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_114 ),
	.cout(Xd_0__inst_mult_28_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_12_q ),
	.datab(!Xd_0__inst_mult_27_13_q ),
	.datac(!Xd_0__inst_mult_27_14_q ),
	.datad(!Xd_0__inst_mult_27_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_114 ),
	.cout(Xd_0__inst_mult_27_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_12_q ),
	.datab(!Xd_0__inst_mult_26_13_q ),
	.datac(!Xd_0__inst_mult_26_14_q ),
	.datad(!Xd_0__inst_mult_26_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_114 ),
	.cout(Xd_0__inst_mult_26_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_12_q ),
	.datab(!Xd_0__inst_mult_25_13_q ),
	.datac(!Xd_0__inst_mult_25_14_q ),
	.datad(!Xd_0__inst_mult_25_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_114 ),
	.cout(Xd_0__inst_mult_25_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_12_q ),
	.datab(!Xd_0__inst_mult_24_13_q ),
	.datac(!Xd_0__inst_mult_24_14_q ),
	.datad(!Xd_0__inst_mult_24_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_114 ),
	.cout(Xd_0__inst_mult_24_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_12_q ),
	.datab(!Xd_0__inst_mult_23_13_q ),
	.datac(!Xd_0__inst_mult_23_14_q ),
	.datad(!Xd_0__inst_mult_23_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_114 ),
	.cout(Xd_0__inst_mult_23_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_12_q ),
	.datab(!Xd_0__inst_mult_22_13_q ),
	.datac(!Xd_0__inst_mult_22_14_q ),
	.datad(!Xd_0__inst_mult_22_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_114 ),
	.cout(Xd_0__inst_mult_22_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_12_q ),
	.datab(!Xd_0__inst_mult_21_13_q ),
	.datac(!Xd_0__inst_mult_21_14_q ),
	.datad(!Xd_0__inst_mult_21_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_114 ),
	.cout(Xd_0__inst_mult_21_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_12_q ),
	.datab(!Xd_0__inst_mult_20_13_q ),
	.datac(!Xd_0__inst_mult_20_14_q ),
	.datad(!Xd_0__inst_mult_20_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_118 ),
	.cout(Xd_0__inst_mult_20_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_12_q ),
	.datab(!Xd_0__inst_mult_19_13_q ),
	.datac(!Xd_0__inst_mult_19_14_q ),
	.datad(!Xd_0__inst_mult_19_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_118 ),
	.cout(Xd_0__inst_mult_19_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_12_q ),
	.datab(!Xd_0__inst_mult_18_13_q ),
	.datac(!Xd_0__inst_mult_18_14_q ),
	.datad(!Xd_0__inst_mult_18_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_118 ),
	.cout(Xd_0__inst_mult_18_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_12_q ),
	.datab(!Xd_0__inst_mult_17_13_q ),
	.datac(!Xd_0__inst_mult_17_14_q ),
	.datad(!Xd_0__inst_mult_17_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_118 ),
	.cout(Xd_0__inst_mult_17_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_12_q ),
	.datab(!Xd_0__inst_mult_16_13_q ),
	.datac(!Xd_0__inst_mult_16_14_q ),
	.datad(!Xd_0__inst_mult_16_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_118 ),
	.cout(Xd_0__inst_mult_16_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_12_q ),
	.datab(!Xd_0__inst_mult_15_13_q ),
	.datac(!Xd_0__inst_mult_15_14_q ),
	.datad(!Xd_0__inst_mult_15_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_118 ),
	.cout(Xd_0__inst_mult_15_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_12_q ),
	.datab(!Xd_0__inst_mult_14_13_q ),
	.datac(!Xd_0__inst_mult_14_14_q ),
	.datad(!Xd_0__inst_mult_14_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_118 ),
	.cout(Xd_0__inst_mult_14_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_12_q ),
	.datab(!Xd_0__inst_mult_13_13_q ),
	.datac(!Xd_0__inst_mult_13_14_q ),
	.datad(!Xd_0__inst_mult_13_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_118 ),
	.cout(Xd_0__inst_mult_13_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_12_q ),
	.datab(!Xd_0__inst_mult_12_13_q ),
	.datac(!Xd_0__inst_mult_12_14_q ),
	.datad(!Xd_0__inst_mult_12_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_118 ),
	.cout(Xd_0__inst_mult_12_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_12_q ),
	.datab(!Xd_0__inst_mult_11_13_q ),
	.datac(!Xd_0__inst_mult_11_14_q ),
	.datad(!Xd_0__inst_mult_11_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_118 ),
	.cout(Xd_0__inst_mult_11_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_12_q ),
	.datab(!Xd_0__inst_mult_10_13_q ),
	.datac(!Xd_0__inst_mult_10_14_q ),
	.datad(!Xd_0__inst_mult_10_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_118 ),
	.cout(Xd_0__inst_mult_10_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_12_q ),
	.datab(!Xd_0__inst_mult_9_13_q ),
	.datac(!Xd_0__inst_mult_9_14_q ),
	.datad(!Xd_0__inst_mult_9_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_118 ),
	.cout(Xd_0__inst_mult_9_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_12_q ),
	.datab(!Xd_0__inst_mult_8_13_q ),
	.datac(!Xd_0__inst_mult_8_14_q ),
	.datad(!Xd_0__inst_mult_8_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_118 ),
	.cout(Xd_0__inst_mult_8_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_12_q ),
	.datab(!Xd_0__inst_mult_7_13_q ),
	.datac(!Xd_0__inst_mult_7_14_q ),
	.datad(!Xd_0__inst_mult_7_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_118 ),
	.cout(Xd_0__inst_mult_7_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_12_q ),
	.datab(!Xd_0__inst_mult_6_13_q ),
	.datac(!Xd_0__inst_mult_6_14_q ),
	.datad(!Xd_0__inst_mult_6_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_118 ),
	.cout(Xd_0__inst_mult_6_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_12_q ),
	.datab(!Xd_0__inst_mult_5_13_q ),
	.datac(!Xd_0__inst_mult_5_14_q ),
	.datad(!Xd_0__inst_mult_5_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_114 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_118 ),
	.cout(Xd_0__inst_mult_5_119 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_12_q ),
	.datab(!Xd_0__inst_mult_4_13_q ),
	.datac(!Xd_0__inst_mult_4_14_q ),
	.datad(!Xd_0__inst_mult_4_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_114 ),
	.cout(Xd_0__inst_mult_4_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_12_q ),
	.datab(!Xd_0__inst_mult_3_13_q ),
	.datac(!Xd_0__inst_mult_3_14_q ),
	.datad(!Xd_0__inst_mult_3_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_114 ),
	.cout(Xd_0__inst_mult_3_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_12_q ),
	.datab(!Xd_0__inst_mult_2_13_q ),
	.datac(!Xd_0__inst_mult_2_14_q ),
	.datad(!Xd_0__inst_mult_2_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_114 ),
	.cout(Xd_0__inst_mult_2_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_12_q ),
	.datab(!Xd_0__inst_mult_1_13_q ),
	.datac(!Xd_0__inst_mult_1_14_q ),
	.datad(!Xd_0__inst_mult_1_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_114 ),
	.cout(Xd_0__inst_mult_1_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_12_q ),
	.datab(!Xd_0__inst_mult_0_13_q ),
	.datac(!Xd_0__inst_mult_0_14_q ),
	.datad(!Xd_0__inst_mult_0_15_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_110 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_114 ),
	.cout(Xd_0__inst_mult_0_115 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_16_q ),
	.datab(!Xd_0__inst_mult_31_17_q ),
	.datac(!Xd_0__inst_mult_31_12_q ),
	.datad(!Xd_0__inst_mult_31_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_119 ),
	.cout(Xd_0__inst_mult_31_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_16_q ),
	.datab(!Xd_0__inst_mult_30_17_q ),
	.datac(!Xd_0__inst_mult_30_12_q ),
	.datad(!Xd_0__inst_mult_30_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_119 ),
	.cout(Xd_0__inst_mult_30_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_16_q ),
	.datab(!Xd_0__inst_mult_29_17_q ),
	.datac(!Xd_0__inst_mult_29_12_q ),
	.datad(!Xd_0__inst_mult_29_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_119 ),
	.cout(Xd_0__inst_mult_29_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_16_q ),
	.datab(!Xd_0__inst_mult_28_17_q ),
	.datac(!Xd_0__inst_mult_28_12_q ),
	.datad(!Xd_0__inst_mult_28_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_119 ),
	.cout(Xd_0__inst_mult_28_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_16_q ),
	.datab(!Xd_0__inst_mult_27_17_q ),
	.datac(!Xd_0__inst_mult_27_12_q ),
	.datad(!Xd_0__inst_mult_27_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_119 ),
	.cout(Xd_0__inst_mult_27_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_16_q ),
	.datab(!Xd_0__inst_mult_26_17_q ),
	.datac(!Xd_0__inst_mult_26_12_q ),
	.datad(!Xd_0__inst_mult_26_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_119 ),
	.cout(Xd_0__inst_mult_26_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_16_q ),
	.datab(!Xd_0__inst_mult_25_17_q ),
	.datac(!Xd_0__inst_mult_25_12_q ),
	.datad(!Xd_0__inst_mult_25_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_119 ),
	.cout(Xd_0__inst_mult_25_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_16_q ),
	.datab(!Xd_0__inst_mult_24_17_q ),
	.datac(!Xd_0__inst_mult_24_12_q ),
	.datad(!Xd_0__inst_mult_24_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_119 ),
	.cout(Xd_0__inst_mult_24_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_16_q ),
	.datab(!Xd_0__inst_mult_23_17_q ),
	.datac(!Xd_0__inst_mult_23_12_q ),
	.datad(!Xd_0__inst_mult_23_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_119 ),
	.cout(Xd_0__inst_mult_23_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_16_q ),
	.datab(!Xd_0__inst_mult_22_17_q ),
	.datac(!Xd_0__inst_mult_22_12_q ),
	.datad(!Xd_0__inst_mult_22_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_119 ),
	.cout(Xd_0__inst_mult_22_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_16_q ),
	.datab(!Xd_0__inst_mult_21_17_q ),
	.datac(!Xd_0__inst_mult_21_12_q ),
	.datad(!Xd_0__inst_mult_21_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_119 ),
	.cout(Xd_0__inst_mult_21_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_16_q ),
	.datab(!Xd_0__inst_mult_20_17_q ),
	.datac(!Xd_0__inst_mult_20_12_q ),
	.datad(!Xd_0__inst_mult_20_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_123 ),
	.cout(Xd_0__inst_mult_20_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_16_q ),
	.datab(!Xd_0__inst_mult_19_17_q ),
	.datac(!Xd_0__inst_mult_19_12_q ),
	.datad(!Xd_0__inst_mult_19_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_123 ),
	.cout(Xd_0__inst_mult_19_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_16_q ),
	.datab(!Xd_0__inst_mult_18_17_q ),
	.datac(!Xd_0__inst_mult_18_12_q ),
	.datad(!Xd_0__inst_mult_18_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_123 ),
	.cout(Xd_0__inst_mult_18_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_16_q ),
	.datab(!Xd_0__inst_mult_17_17_q ),
	.datac(!Xd_0__inst_mult_17_12_q ),
	.datad(!Xd_0__inst_mult_17_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_123 ),
	.cout(Xd_0__inst_mult_17_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_16_q ),
	.datab(!Xd_0__inst_mult_16_17_q ),
	.datac(!Xd_0__inst_mult_16_12_q ),
	.datad(!Xd_0__inst_mult_16_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_123 ),
	.cout(Xd_0__inst_mult_16_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_16_q ),
	.datab(!Xd_0__inst_mult_15_17_q ),
	.datac(!Xd_0__inst_mult_15_12_q ),
	.datad(!Xd_0__inst_mult_15_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_123 ),
	.cout(Xd_0__inst_mult_15_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_16_q ),
	.datab(!Xd_0__inst_mult_14_17_q ),
	.datac(!Xd_0__inst_mult_14_12_q ),
	.datad(!Xd_0__inst_mult_14_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_123 ),
	.cout(Xd_0__inst_mult_14_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_16_q ),
	.datab(!Xd_0__inst_mult_13_17_q ),
	.datac(!Xd_0__inst_mult_13_12_q ),
	.datad(!Xd_0__inst_mult_13_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_123 ),
	.cout(Xd_0__inst_mult_13_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_16_q ),
	.datab(!Xd_0__inst_mult_12_17_q ),
	.datac(!Xd_0__inst_mult_12_12_q ),
	.datad(!Xd_0__inst_mult_12_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_123 ),
	.cout(Xd_0__inst_mult_12_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_16_q ),
	.datab(!Xd_0__inst_mult_11_17_q ),
	.datac(!Xd_0__inst_mult_11_12_q ),
	.datad(!Xd_0__inst_mult_11_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_123 ),
	.cout(Xd_0__inst_mult_11_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_16_q ),
	.datab(!Xd_0__inst_mult_10_17_q ),
	.datac(!Xd_0__inst_mult_10_12_q ),
	.datad(!Xd_0__inst_mult_10_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_123 ),
	.cout(Xd_0__inst_mult_10_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_16_q ),
	.datab(!Xd_0__inst_mult_9_17_q ),
	.datac(!Xd_0__inst_mult_9_12_q ),
	.datad(!Xd_0__inst_mult_9_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_123 ),
	.cout(Xd_0__inst_mult_9_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_16_q ),
	.datab(!Xd_0__inst_mult_8_17_q ),
	.datac(!Xd_0__inst_mult_8_12_q ),
	.datad(!Xd_0__inst_mult_8_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_123 ),
	.cout(Xd_0__inst_mult_8_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_16_q ),
	.datab(!Xd_0__inst_mult_7_17_q ),
	.datac(!Xd_0__inst_mult_7_12_q ),
	.datad(!Xd_0__inst_mult_7_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_123 ),
	.cout(Xd_0__inst_mult_7_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_16_q ),
	.datab(!Xd_0__inst_mult_6_17_q ),
	.datac(!Xd_0__inst_mult_6_12_q ),
	.datad(!Xd_0__inst_mult_6_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_123 ),
	.cout(Xd_0__inst_mult_6_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_16_q ),
	.datab(!Xd_0__inst_mult_5_17_q ),
	.datac(!Xd_0__inst_mult_5_12_q ),
	.datad(!Xd_0__inst_mult_5_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_119 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_123 ),
	.cout(Xd_0__inst_mult_5_124 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_16_q ),
	.datab(!Xd_0__inst_mult_4_17_q ),
	.datac(!Xd_0__inst_mult_4_12_q ),
	.datad(!Xd_0__inst_mult_4_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_119 ),
	.cout(Xd_0__inst_mult_4_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_16_q ),
	.datab(!Xd_0__inst_mult_3_17_q ),
	.datac(!Xd_0__inst_mult_3_12_q ),
	.datad(!Xd_0__inst_mult_3_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_119 ),
	.cout(Xd_0__inst_mult_3_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_16_q ),
	.datab(!Xd_0__inst_mult_2_17_q ),
	.datac(!Xd_0__inst_mult_2_12_q ),
	.datad(!Xd_0__inst_mult_2_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_119 ),
	.cout(Xd_0__inst_mult_2_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_16_q ),
	.datab(!Xd_0__inst_mult_1_17_q ),
	.datac(!Xd_0__inst_mult_1_12_q ),
	.datad(!Xd_0__inst_mult_1_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_119 ),
	.cout(Xd_0__inst_mult_1_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_42 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_16_q ),
	.datab(!Xd_0__inst_mult_0_17_q ),
	.datac(!Xd_0__inst_mult_0_12_q ),
	.datad(!Xd_0__inst_mult_0_13_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_115 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_119 ),
	.cout(Xd_0__inst_mult_0_120 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_18_q ),
	.datab(!Xd_0__inst_mult_31_19_q ),
	.datac(!Xd_0__inst_mult_31_16_q ),
	.datad(!Xd_0__inst_mult_31_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_124 ),
	.cout(Xd_0__inst_mult_31_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_18_q ),
	.datab(!Xd_0__inst_mult_30_19_q ),
	.datac(!Xd_0__inst_mult_30_16_q ),
	.datad(!Xd_0__inst_mult_30_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_124 ),
	.cout(Xd_0__inst_mult_30_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_18_q ),
	.datab(!Xd_0__inst_mult_29_19_q ),
	.datac(!Xd_0__inst_mult_29_16_q ),
	.datad(!Xd_0__inst_mult_29_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_124 ),
	.cout(Xd_0__inst_mult_29_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_18_q ),
	.datab(!Xd_0__inst_mult_28_19_q ),
	.datac(!Xd_0__inst_mult_28_16_q ),
	.datad(!Xd_0__inst_mult_28_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_124 ),
	.cout(Xd_0__inst_mult_28_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_18_q ),
	.datab(!Xd_0__inst_mult_27_19_q ),
	.datac(!Xd_0__inst_mult_27_16_q ),
	.datad(!Xd_0__inst_mult_27_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_124 ),
	.cout(Xd_0__inst_mult_27_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_18_q ),
	.datab(!Xd_0__inst_mult_26_19_q ),
	.datac(!Xd_0__inst_mult_26_16_q ),
	.datad(!Xd_0__inst_mult_26_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_124 ),
	.cout(Xd_0__inst_mult_26_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_18_q ),
	.datab(!Xd_0__inst_mult_25_19_q ),
	.datac(!Xd_0__inst_mult_25_16_q ),
	.datad(!Xd_0__inst_mult_25_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_124 ),
	.cout(Xd_0__inst_mult_25_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_18_q ),
	.datab(!Xd_0__inst_mult_24_19_q ),
	.datac(!Xd_0__inst_mult_24_16_q ),
	.datad(!Xd_0__inst_mult_24_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_124 ),
	.cout(Xd_0__inst_mult_24_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_18_q ),
	.datab(!Xd_0__inst_mult_23_19_q ),
	.datac(!Xd_0__inst_mult_23_16_q ),
	.datad(!Xd_0__inst_mult_23_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_124 ),
	.cout(Xd_0__inst_mult_23_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_18_q ),
	.datab(!Xd_0__inst_mult_22_19_q ),
	.datac(!Xd_0__inst_mult_22_16_q ),
	.datad(!Xd_0__inst_mult_22_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_124 ),
	.cout(Xd_0__inst_mult_22_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_18_q ),
	.datab(!Xd_0__inst_mult_21_19_q ),
	.datac(!Xd_0__inst_mult_21_16_q ),
	.datad(!Xd_0__inst_mult_21_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_124 ),
	.cout(Xd_0__inst_mult_21_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_18_q ),
	.datab(!Xd_0__inst_mult_20_19_q ),
	.datac(!Xd_0__inst_mult_20_16_q ),
	.datad(!Xd_0__inst_mult_20_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_128 ),
	.cout(Xd_0__inst_mult_20_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_18_q ),
	.datab(!Xd_0__inst_mult_19_19_q ),
	.datac(!Xd_0__inst_mult_19_16_q ),
	.datad(!Xd_0__inst_mult_19_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_128 ),
	.cout(Xd_0__inst_mult_19_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_18_q ),
	.datab(!Xd_0__inst_mult_18_19_q ),
	.datac(!Xd_0__inst_mult_18_16_q ),
	.datad(!Xd_0__inst_mult_18_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_128 ),
	.cout(Xd_0__inst_mult_18_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_18_q ),
	.datab(!Xd_0__inst_mult_17_19_q ),
	.datac(!Xd_0__inst_mult_17_16_q ),
	.datad(!Xd_0__inst_mult_17_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_128 ),
	.cout(Xd_0__inst_mult_17_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_18_q ),
	.datab(!Xd_0__inst_mult_16_19_q ),
	.datac(!Xd_0__inst_mult_16_16_q ),
	.datad(!Xd_0__inst_mult_16_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_128 ),
	.cout(Xd_0__inst_mult_16_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_18_q ),
	.datab(!Xd_0__inst_mult_15_19_q ),
	.datac(!Xd_0__inst_mult_15_16_q ),
	.datad(!Xd_0__inst_mult_15_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_128 ),
	.cout(Xd_0__inst_mult_15_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_18_q ),
	.datab(!Xd_0__inst_mult_14_19_q ),
	.datac(!Xd_0__inst_mult_14_16_q ),
	.datad(!Xd_0__inst_mult_14_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_128 ),
	.cout(Xd_0__inst_mult_14_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_18_q ),
	.datab(!Xd_0__inst_mult_13_19_q ),
	.datac(!Xd_0__inst_mult_13_16_q ),
	.datad(!Xd_0__inst_mult_13_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_128 ),
	.cout(Xd_0__inst_mult_13_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_18_q ),
	.datab(!Xd_0__inst_mult_12_19_q ),
	.datac(!Xd_0__inst_mult_12_16_q ),
	.datad(!Xd_0__inst_mult_12_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_128 ),
	.cout(Xd_0__inst_mult_12_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_18_q ),
	.datab(!Xd_0__inst_mult_11_19_q ),
	.datac(!Xd_0__inst_mult_11_16_q ),
	.datad(!Xd_0__inst_mult_11_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_128 ),
	.cout(Xd_0__inst_mult_11_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_18_q ),
	.datab(!Xd_0__inst_mult_10_19_q ),
	.datac(!Xd_0__inst_mult_10_16_q ),
	.datad(!Xd_0__inst_mult_10_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_128 ),
	.cout(Xd_0__inst_mult_10_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_18_q ),
	.datab(!Xd_0__inst_mult_9_19_q ),
	.datac(!Xd_0__inst_mult_9_16_q ),
	.datad(!Xd_0__inst_mult_9_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_128 ),
	.cout(Xd_0__inst_mult_9_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_18_q ),
	.datab(!Xd_0__inst_mult_8_19_q ),
	.datac(!Xd_0__inst_mult_8_16_q ),
	.datad(!Xd_0__inst_mult_8_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_128 ),
	.cout(Xd_0__inst_mult_8_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_18_q ),
	.datab(!Xd_0__inst_mult_7_19_q ),
	.datac(!Xd_0__inst_mult_7_16_q ),
	.datad(!Xd_0__inst_mult_7_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_128 ),
	.cout(Xd_0__inst_mult_7_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_18_q ),
	.datab(!Xd_0__inst_mult_6_19_q ),
	.datac(!Xd_0__inst_mult_6_16_q ),
	.datad(!Xd_0__inst_mult_6_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_128 ),
	.cout(Xd_0__inst_mult_6_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_18_q ),
	.datab(!Xd_0__inst_mult_5_19_q ),
	.datac(!Xd_0__inst_mult_5_16_q ),
	.datad(!Xd_0__inst_mult_5_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_124 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_128 ),
	.cout(Xd_0__inst_mult_5_129 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_18_q ),
	.datab(!Xd_0__inst_mult_4_19_q ),
	.datac(!Xd_0__inst_mult_4_16_q ),
	.datad(!Xd_0__inst_mult_4_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_124 ),
	.cout(Xd_0__inst_mult_4_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_18_q ),
	.datab(!Xd_0__inst_mult_3_19_q ),
	.datac(!Xd_0__inst_mult_3_16_q ),
	.datad(!Xd_0__inst_mult_3_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_124 ),
	.cout(Xd_0__inst_mult_3_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_18_q ),
	.datab(!Xd_0__inst_mult_2_19_q ),
	.datac(!Xd_0__inst_mult_2_16_q ),
	.datad(!Xd_0__inst_mult_2_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_124 ),
	.cout(Xd_0__inst_mult_2_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_18_q ),
	.datab(!Xd_0__inst_mult_1_19_q ),
	.datac(!Xd_0__inst_mult_1_16_q ),
	.datad(!Xd_0__inst_mult_1_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_124 ),
	.cout(Xd_0__inst_mult_1_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_43 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_18_q ),
	.datab(!Xd_0__inst_mult_0_19_q ),
	.datac(!Xd_0__inst_mult_0_16_q ),
	.datad(!Xd_0__inst_mult_0_17_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_120 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_124 ),
	.cout(Xd_0__inst_mult_0_125 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_20_q ),
	.datab(!Xd_0__inst_mult_31_21_q ),
	.datac(!Xd_0__inst_mult_31_18_q ),
	.datad(!Xd_0__inst_mult_31_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_129 ),
	.cout(Xd_0__inst_mult_31_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_20_q ),
	.datab(!Xd_0__inst_mult_30_21_q ),
	.datac(!Xd_0__inst_mult_30_18_q ),
	.datad(!Xd_0__inst_mult_30_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_129 ),
	.cout(Xd_0__inst_mult_30_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_20_q ),
	.datab(!Xd_0__inst_mult_29_21_q ),
	.datac(!Xd_0__inst_mult_29_18_q ),
	.datad(!Xd_0__inst_mult_29_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_129 ),
	.cout(Xd_0__inst_mult_29_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_20_q ),
	.datab(!Xd_0__inst_mult_28_21_q ),
	.datac(!Xd_0__inst_mult_28_18_q ),
	.datad(!Xd_0__inst_mult_28_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_129 ),
	.cout(Xd_0__inst_mult_28_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_20_q ),
	.datab(!Xd_0__inst_mult_27_21_q ),
	.datac(!Xd_0__inst_mult_27_18_q ),
	.datad(!Xd_0__inst_mult_27_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_129 ),
	.cout(Xd_0__inst_mult_27_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_20_q ),
	.datab(!Xd_0__inst_mult_26_21_q ),
	.datac(!Xd_0__inst_mult_26_18_q ),
	.datad(!Xd_0__inst_mult_26_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_129 ),
	.cout(Xd_0__inst_mult_26_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_20_q ),
	.datab(!Xd_0__inst_mult_25_21_q ),
	.datac(!Xd_0__inst_mult_25_18_q ),
	.datad(!Xd_0__inst_mult_25_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_129 ),
	.cout(Xd_0__inst_mult_25_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_20_q ),
	.datab(!Xd_0__inst_mult_24_21_q ),
	.datac(!Xd_0__inst_mult_24_18_q ),
	.datad(!Xd_0__inst_mult_24_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_129 ),
	.cout(Xd_0__inst_mult_24_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_20_q ),
	.datab(!Xd_0__inst_mult_23_21_q ),
	.datac(!Xd_0__inst_mult_23_18_q ),
	.datad(!Xd_0__inst_mult_23_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_129 ),
	.cout(Xd_0__inst_mult_23_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_20_q ),
	.datab(!Xd_0__inst_mult_22_21_q ),
	.datac(!Xd_0__inst_mult_22_18_q ),
	.datad(!Xd_0__inst_mult_22_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_129 ),
	.cout(Xd_0__inst_mult_22_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_20_q ),
	.datab(!Xd_0__inst_mult_21_21_q ),
	.datac(!Xd_0__inst_mult_21_18_q ),
	.datad(!Xd_0__inst_mult_21_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_129 ),
	.cout(Xd_0__inst_mult_21_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_20_q ),
	.datab(!Xd_0__inst_mult_20_21_q ),
	.datac(!Xd_0__inst_mult_20_18_q ),
	.datad(!Xd_0__inst_mult_20_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_133 ),
	.cout(Xd_0__inst_mult_20_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_20_q ),
	.datab(!Xd_0__inst_mult_19_21_q ),
	.datac(!Xd_0__inst_mult_19_18_q ),
	.datad(!Xd_0__inst_mult_19_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_133 ),
	.cout(Xd_0__inst_mult_19_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_20_q ),
	.datab(!Xd_0__inst_mult_18_21_q ),
	.datac(!Xd_0__inst_mult_18_18_q ),
	.datad(!Xd_0__inst_mult_18_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_133 ),
	.cout(Xd_0__inst_mult_18_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_20_q ),
	.datab(!Xd_0__inst_mult_17_21_q ),
	.datac(!Xd_0__inst_mult_17_18_q ),
	.datad(!Xd_0__inst_mult_17_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_133 ),
	.cout(Xd_0__inst_mult_17_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_20_q ),
	.datab(!Xd_0__inst_mult_16_21_q ),
	.datac(!Xd_0__inst_mult_16_18_q ),
	.datad(!Xd_0__inst_mult_16_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_133 ),
	.cout(Xd_0__inst_mult_16_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_20_q ),
	.datab(!Xd_0__inst_mult_15_21_q ),
	.datac(!Xd_0__inst_mult_15_18_q ),
	.datad(!Xd_0__inst_mult_15_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_133 ),
	.cout(Xd_0__inst_mult_15_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_20_q ),
	.datab(!Xd_0__inst_mult_14_21_q ),
	.datac(!Xd_0__inst_mult_14_18_q ),
	.datad(!Xd_0__inst_mult_14_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_133 ),
	.cout(Xd_0__inst_mult_14_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_20_q ),
	.datab(!Xd_0__inst_mult_13_21_q ),
	.datac(!Xd_0__inst_mult_13_18_q ),
	.datad(!Xd_0__inst_mult_13_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_133 ),
	.cout(Xd_0__inst_mult_13_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_20_q ),
	.datab(!Xd_0__inst_mult_12_21_q ),
	.datac(!Xd_0__inst_mult_12_18_q ),
	.datad(!Xd_0__inst_mult_12_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_133 ),
	.cout(Xd_0__inst_mult_12_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_20_q ),
	.datab(!Xd_0__inst_mult_11_21_q ),
	.datac(!Xd_0__inst_mult_11_18_q ),
	.datad(!Xd_0__inst_mult_11_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_133 ),
	.cout(Xd_0__inst_mult_11_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_20_q ),
	.datab(!Xd_0__inst_mult_10_21_q ),
	.datac(!Xd_0__inst_mult_10_18_q ),
	.datad(!Xd_0__inst_mult_10_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_133 ),
	.cout(Xd_0__inst_mult_10_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_20_q ),
	.datab(!Xd_0__inst_mult_9_21_q ),
	.datac(!Xd_0__inst_mult_9_18_q ),
	.datad(!Xd_0__inst_mult_9_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_133 ),
	.cout(Xd_0__inst_mult_9_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_20_q ),
	.datab(!Xd_0__inst_mult_8_21_q ),
	.datac(!Xd_0__inst_mult_8_18_q ),
	.datad(!Xd_0__inst_mult_8_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_133 ),
	.cout(Xd_0__inst_mult_8_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_20_q ),
	.datab(!Xd_0__inst_mult_7_21_q ),
	.datac(!Xd_0__inst_mult_7_18_q ),
	.datad(!Xd_0__inst_mult_7_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_133 ),
	.cout(Xd_0__inst_mult_7_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_20_q ),
	.datab(!Xd_0__inst_mult_6_21_q ),
	.datac(!Xd_0__inst_mult_6_18_q ),
	.datad(!Xd_0__inst_mult_6_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_133 ),
	.cout(Xd_0__inst_mult_6_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_20_q ),
	.datab(!Xd_0__inst_mult_5_21_q ),
	.datac(!Xd_0__inst_mult_5_18_q ),
	.datad(!Xd_0__inst_mult_5_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_129 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_133 ),
	.cout(Xd_0__inst_mult_5_134 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_20_q ),
	.datab(!Xd_0__inst_mult_4_21_q ),
	.datac(!Xd_0__inst_mult_4_18_q ),
	.datad(!Xd_0__inst_mult_4_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_129 ),
	.cout(Xd_0__inst_mult_4_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_20_q ),
	.datab(!Xd_0__inst_mult_3_21_q ),
	.datac(!Xd_0__inst_mult_3_18_q ),
	.datad(!Xd_0__inst_mult_3_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_129 ),
	.cout(Xd_0__inst_mult_3_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_20_q ),
	.datab(!Xd_0__inst_mult_2_21_q ),
	.datac(!Xd_0__inst_mult_2_18_q ),
	.datad(!Xd_0__inst_mult_2_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_129 ),
	.cout(Xd_0__inst_mult_2_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_20_q ),
	.datab(!Xd_0__inst_mult_1_21_q ),
	.datac(!Xd_0__inst_mult_1_18_q ),
	.datad(!Xd_0__inst_mult_1_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_129 ),
	.cout(Xd_0__inst_mult_1_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_44 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_20_q ),
	.datab(!Xd_0__inst_mult_0_21_q ),
	.datac(!Xd_0__inst_mult_0_18_q ),
	.datad(!Xd_0__inst_mult_0_19_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_125 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_129 ),
	.cout(Xd_0__inst_mult_0_130 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_20_q ),
	.datab(!Xd_0__inst_mult_31_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_20_q ),
	.datab(!Xd_0__inst_mult_30_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_20_q ),
	.datab(!Xd_0__inst_mult_29_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_20_q ),
	.datab(!Xd_0__inst_mult_28_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_20_q ),
	.datab(!Xd_0__inst_mult_27_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_20_q ),
	.datab(!Xd_0__inst_mult_26_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_20_q ),
	.datab(!Xd_0__inst_mult_25_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_20_q ),
	.datab(!Xd_0__inst_mult_24_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_20_q ),
	.datab(!Xd_0__inst_mult_23_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_20_q ),
	.datab(!Xd_0__inst_mult_22_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_20_q ),
	.datab(!Xd_0__inst_mult_21_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_20_q ),
	.datab(!Xd_0__inst_mult_20_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_20_q ),
	.datab(!Xd_0__inst_mult_19_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_20_q ),
	.datab(!Xd_0__inst_mult_18_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_20_q ),
	.datab(!Xd_0__inst_mult_17_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_20_q ),
	.datab(!Xd_0__inst_mult_16_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_20_q ),
	.datab(!Xd_0__inst_mult_15_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_20_q ),
	.datab(!Xd_0__inst_mult_14_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_20_q ),
	.datab(!Xd_0__inst_mult_13_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_20_q ),
	.datab(!Xd_0__inst_mult_12_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_20_q ),
	.datab(!Xd_0__inst_mult_11_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_20_q ),
	.datab(!Xd_0__inst_mult_10_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_20_q ),
	.datab(!Xd_0__inst_mult_9_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_20_q ),
	.datab(!Xd_0__inst_mult_8_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_20_q ),
	.datab(!Xd_0__inst_mult_7_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_20_q ),
	.datab(!Xd_0__inst_mult_6_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_46 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_20_q ),
	.datab(!Xd_0__inst_mult_5_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_134 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_138 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_20_q ),
	.datab(!Xd_0__inst_mult_4_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_20_q ),
	.datab(!Xd_0__inst_mult_3_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_20_q ),
	.datab(!Xd_0__inst_mult_2_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_20_q ),
	.datab(!Xd_0__inst_mult_1_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_45 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_20_q ),
	.datab(!Xd_0__inst_mult_0_21_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_130 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_134 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_41 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[247]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_41_sumout ),
	.cout(Xd_0__inst_i21_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_31_46 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[248]),
	.datac(!din_a[249]),
	.datad(!din_b[249]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_139 ),
	.cout(Xd_0__inst_mult_31_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_30_46 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[240]),
	.datac(!din_a[241]),
	.datad(!din_b[241]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_139 ),
	.cout(Xd_0__inst_mult_30_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_47 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[45]),
	.datac(!din_a[44]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_143 ),
	.cout(Xd_0__inst_mult_5_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_46 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[231]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_46_sumout ),
	.cout(Xd_0__inst_i21_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_51 (
// Equation(s):

	.dataa(!din_a[239]),
	.datab(!din_b[239]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_51_sumout ),
	.cout(Xd_0__inst_i21_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_29_46 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[232]),
	.datac(!din_a[233]),
	.datad(!din_b[233]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_139 ),
	.cout(Xd_0__inst_mult_29_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_28_46 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[224]),
	.datac(!din_a[225]),
	.datad(!din_b[225]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_139 ),
	.cout(Xd_0__inst_mult_28_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_47 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[53]),
	.datac(!din_a[52]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_143 ),
	.cout(Xd_0__inst_mult_6_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_56 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_56_sumout ),
	.cout(Xd_0__inst_i21_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_61 (
// Equation(s):

	.dataa(!din_a[215]),
	.datab(!din_b[215]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_61_sumout ),
	.cout(Xd_0__inst_i21_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_27_46 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[216]),
	.datac(!din_a[217]),
	.datad(!din_b[217]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_139 ),
	.cout(Xd_0__inst_mult_27_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_26_46 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[208]),
	.datac(!din_a[209]),
	.datad(!din_b[209]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_139 ),
	.cout(Xd_0__inst_mult_26_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_47 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[61]),
	.datac(!din_a[60]),
	.datad(!din_b[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_143 ),
	.cout(Xd_0__inst_mult_7_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_66 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[199]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_66_sumout ),
	.cout(Xd_0__inst_i21_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_71 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[207]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_71_sumout ),
	.cout(Xd_0__inst_i21_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_25_46 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[200]),
	.datac(!din_a[201]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_139 ),
	.cout(Xd_0__inst_mult_25_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_24_46 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[192]),
	.datac(!din_a[193]),
	.datad(!din_b[193]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_139 ),
	.cout(Xd_0__inst_mult_24_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_47 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[69]),
	.datac(!din_a[68]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_143 ),
	.cout(Xd_0__inst_mult_8_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_76 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[183]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_76_sumout ),
	.cout(Xd_0__inst_i21_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_23_46 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[184]),
	.datac(!din_a[185]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_139 ),
	.cout(Xd_0__inst_mult_23_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_22_46 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[176]),
	.datac(!din_a[177]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_139 ),
	.cout(Xd_0__inst_mult_22_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_47 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[77]),
	.datac(!din_a[76]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_143 ),
	.cout(Xd_0__inst_mult_9_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_81 (
// Equation(s):

	.dataa(!din_a[167]),
	.datab(!din_b[167]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_81_sumout ),
	.cout(Xd_0__inst_i21_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_86 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[175]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_86_sumout ),
	.cout(Xd_0__inst_i21_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_21_46 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[168]),
	.datac(!din_a[169]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_139 ),
	.cout(Xd_0__inst_mult_21_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_20_47 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[160]),
	.datac(!din_a[161]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_143 ),
	.cout(Xd_0__inst_mult_20_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_48 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[165]),
	.datac(!din_a[164]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_148 ),
	.cout(Xd_0__inst_mult_20_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_19_47 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[152]),
	.datac(!din_a[153]),
	.datad(!din_b[153]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_143 ),
	.cout(Xd_0__inst_mult_19_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_18_47 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[144]),
	.datac(!din_a[145]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_143 ),
	.cout(Xd_0__inst_mult_18_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_48 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[157]),
	.datac(!din_a[156]),
	.datad(!din_b[155]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_148 ),
	.cout(Xd_0__inst_mult_19_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_91 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[135]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_91_sumout ),
	.cout(Xd_0__inst_i21_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_96 (
// Equation(s):

	.dataa(!din_a[143]),
	.datab(!din_b[143]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_96_sumout ),
	.cout(Xd_0__inst_i21_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_17_47 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[136]),
	.datac(!din_a[137]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_143 ),
	.cout(Xd_0__inst_mult_17_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_16_47 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[128]),
	.datac(!din_a[129]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_143 ),
	.cout(Xd_0__inst_mult_16_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_47 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[93]),
	.datac(!din_a[92]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_143 ),
	.cout(Xd_0__inst_mult_11_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_101 (
// Equation(s):

	.dataa(!din_a[119]),
	.datab(!din_b[119]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_101_sumout ),
	.cout(Xd_0__inst_i21_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_15_47 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[120]),
	.datac(!din_a[121]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_143 ),
	.cout(Xd_0__inst_mult_15_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_14_47 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[112]),
	.datac(!din_a[113]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_143 ),
	.cout(Xd_0__inst_mult_14_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_48 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[149]),
	.datac(!din_a[148]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_148 ),
	.cout(Xd_0__inst_mult_18_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_106 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_106_sumout ),
	.cout(Xd_0__inst_i21_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_111 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[111]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_111_sumout ),
	.cout(Xd_0__inst_i21_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_13_47 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[104]),
	.datac(!din_a[105]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_143 ),
	.cout(Xd_0__inst_mult_13_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_12_47 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[96]),
	.datac(!din_a[97]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_143 ),
	.cout(Xd_0__inst_mult_12_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_48 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[141]),
	.datac(!din_a[140]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_148 ),
	.cout(Xd_0__inst_mult_17_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_116 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[87]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_116_sumout ),
	.cout(Xd_0__inst_i21_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_11_48 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[88]),
	.datac(!din_a[89]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_148 ),
	.cout(Xd_0__inst_mult_11_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_10_47 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[80]),
	.datac(!din_a[81]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_143 ),
	.cout(Xd_0__inst_mult_10_144 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_48 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[133]),
	.datac(!din_a[132]),
	.datad(!din_b[131]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_148 ),
	.cout(Xd_0__inst_mult_16_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_121 (
// Equation(s):

	.dataa(!din_a[71]),
	.datab(!din_b[71]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_127 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_121_sumout ),
	.cout(Xd_0__inst_i21_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_126 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_126_sumout ),
	.cout(Xd_0__inst_i21_127 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_9_48 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(!din_a[73]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_148 ),
	.cout(Xd_0__inst_mult_9_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_8_48 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[64]),
	.datac(!din_a[65]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_148 ),
	.cout(Xd_0__inst_mult_8_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_48 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[85]),
	.datac(!din_a[84]),
	.datad(!din_b[83]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_148 ),
	.cout(Xd_0__inst_mult_10_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_131 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_137 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_131_sumout ),
	.cout(Xd_0__inst_i21_132 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_7_48 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[56]),
	.datac(!din_a[57]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_148 ),
	.cout(Xd_0__inst_mult_7_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_6_48 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(!din_a[49]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_148 ),
	.cout(Xd_0__inst_mult_6_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_48 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[125]),
	.datac(!din_a[124]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_148 ),
	.cout(Xd_0__inst_mult_15_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_136 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[39]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_142 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_136_sumout ),
	.cout(Xd_0__inst_i21_137 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_141 (
// Equation(s):

	.dataa(!din_a[47]),
	.datab(!din_b[47]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_147 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_141_sumout ),
	.cout(Xd_0__inst_i21_142 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_5_48 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[40]),
	.datac(!din_a[41]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_154 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_148 ),
	.cout(Xd_0__inst_mult_5_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_4_46 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[32]),
	.datac(!din_a[33]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_139 ),
	.cout(Xd_0__inst_mult_4_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_48 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[117]),
	.datac(!din_a[116]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_148 ),
	.cout(Xd_0__inst_mult_14_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_146 (
// Equation(s):

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_146_sumout ),
	.cout(Xd_0__inst_i21_147 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_3_46 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[24]),
	.datac(!din_a[25]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_139 ),
	.cout(Xd_0__inst_mult_3_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_2_46 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[16]),
	.datac(!din_a[17]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_139 ),
	.cout(Xd_0__inst_mult_2_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_48 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[109]),
	.datac(!din_a[108]),
	.datad(!din_b[107]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_148 ),
	.cout(Xd_0__inst_mult_13_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_151 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_157 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_151_sumout ),
	.cout(Xd_0__inst_i21_152 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i21_156 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[15]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i21_156_sumout ),
	.cout(Xd_0__inst_i21_157 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_1_46 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[8]),
	.datac(!din_a[9]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_139 ),
	.cout(Xd_0__inst_mult_1_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_0_46 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(!din_a[1]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_145 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_139 ),
	.cout(Xd_0__inst_mult_0_140 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_48 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[101]),
	.datac(!din_a[100]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_169 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_148 ),
	.cout(Xd_0__inst_mult_12_149 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_47 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[248]),
	.datac(!din_a[248]),
	.datad(!din_b[249]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_144 ),
	.cout(Xd_0__inst_mult_31_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_47 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[240]),
	.datac(!din_a[240]),
	.datad(!din_b[241]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_144 ),
	.cout(Xd_0__inst_mult_30_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_47 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[232]),
	.datac(!din_a[232]),
	.datad(!din_b[233]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_144 ),
	.cout(Xd_0__inst_mult_29_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_47 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[224]),
	.datac(!din_a[224]),
	.datad(!din_b[225]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_144 ),
	.cout(Xd_0__inst_mult_28_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_47 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[216]),
	.datac(!din_a[216]),
	.datad(!din_b[217]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_144 ),
	.cout(Xd_0__inst_mult_27_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_47 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[208]),
	.datac(!din_a[208]),
	.datad(!din_b[209]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_144 ),
	.cout(Xd_0__inst_mult_26_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_47 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[200]),
	.datac(!din_a[200]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_144 ),
	.cout(Xd_0__inst_mult_25_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_47 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[192]),
	.datac(!din_a[192]),
	.datad(!din_b[193]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_144 ),
	.cout(Xd_0__inst_mult_24_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_47 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[184]),
	.datac(!din_a[184]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_144 ),
	.cout(Xd_0__inst_mult_23_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_47 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[176]),
	.datac(!din_a[176]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_144 ),
	.cout(Xd_0__inst_mult_22_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_47 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[168]),
	.datac(!din_a[168]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_144 ),
	.cout(Xd_0__inst_mult_21_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_49 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[160]),
	.datac(!din_a[160]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_153 ),
	.cout(Xd_0__inst_mult_20_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_49 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[152]),
	.datac(!din_a[152]),
	.datad(!din_b[153]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_153 ),
	.cout(Xd_0__inst_mult_19_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_49 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[144]),
	.datac(!din_a[144]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_153 ),
	.cout(Xd_0__inst_mult_18_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_49 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[136]),
	.datac(!din_a[136]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_153 ),
	.cout(Xd_0__inst_mult_17_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_49 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[128]),
	.datac(!din_a[128]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_153 ),
	.cout(Xd_0__inst_mult_16_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_49 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[120]),
	.datac(!din_a[120]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_153 ),
	.cout(Xd_0__inst_mult_15_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_49 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[112]),
	.datac(!din_a[112]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_153 ),
	.cout(Xd_0__inst_mult_14_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_49 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[104]),
	.datac(!din_a[104]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_153 ),
	.cout(Xd_0__inst_mult_13_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_49 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[96]),
	.datac(!din_a[96]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_153 ),
	.cout(Xd_0__inst_mult_12_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_49 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[88]),
	.datac(!din_a[88]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_153 ),
	.cout(Xd_0__inst_mult_11_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_49 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[80]),
	.datac(!din_a[80]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_153 ),
	.cout(Xd_0__inst_mult_10_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_49 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[72]),
	.datac(!din_a[72]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_153 ),
	.cout(Xd_0__inst_mult_9_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_49 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[64]),
	.datac(!din_a[64]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_153 ),
	.cout(Xd_0__inst_mult_8_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_49 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[56]),
	.datac(!din_a[56]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_153 ),
	.cout(Xd_0__inst_mult_7_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_49 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[48]),
	.datac(!din_a[48]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_153 ),
	.cout(Xd_0__inst_mult_6_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_49 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[40]),
	.datac(!din_a[40]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_153 ),
	.cout(Xd_0__inst_mult_5_154 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_47 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[32]),
	.datac(!din_a[32]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_144 ),
	.cout(Xd_0__inst_mult_4_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_47 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[24]),
	.datac(!din_a[24]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_144 ),
	.cout(Xd_0__inst_mult_3_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_47 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[16]),
	.datac(!din_a[16]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_144 ),
	.cout(Xd_0__inst_mult_2_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_47 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[8]),
	.datac(!din_a[8]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_144 ),
	.cout(Xd_0__inst_mult_1_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_47 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[0]),
	.datac(!din_a[0]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_144 ),
	.cout(Xd_0__inst_mult_0_145 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_48 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[248]),
	.datac(!din_a[248]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_149 ),
	.cout(Xd_0__inst_mult_31_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_48 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[240]),
	.datac(!din_a[240]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_149 ),
	.cout(Xd_0__inst_mult_30_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_48 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[232]),
	.datac(!din_a[232]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_149 ),
	.cout(Xd_0__inst_mult_29_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_48 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[224]),
	.datac(!din_a[224]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_149 ),
	.cout(Xd_0__inst_mult_28_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_48 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[216]),
	.datac(!din_a[216]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_149 ),
	.cout(Xd_0__inst_mult_27_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_48 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[208]),
	.datac(!din_a[208]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_149 ),
	.cout(Xd_0__inst_mult_26_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_48 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[200]),
	.datac(!din_a[200]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_149 ),
	.cout(Xd_0__inst_mult_25_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_48 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[192]),
	.datac(!din_a[192]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_149 ),
	.cout(Xd_0__inst_mult_24_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_48 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[184]),
	.datac(!din_a[184]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_149 ),
	.cout(Xd_0__inst_mult_23_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_48 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[176]),
	.datac(!din_a[176]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_149 ),
	.cout(Xd_0__inst_mult_22_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_48 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[168]),
	.datac(!din_a[168]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_149 ),
	.cout(Xd_0__inst_mult_21_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_50 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[160]),
	.datac(!din_a[160]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_158 ),
	.cout(Xd_0__inst_mult_20_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_50 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[152]),
	.datac(!din_a[152]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_158 ),
	.cout(Xd_0__inst_mult_19_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_50 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[144]),
	.datac(!din_a[144]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_158 ),
	.cout(Xd_0__inst_mult_18_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_50 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[136]),
	.datac(!din_a[136]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_158 ),
	.cout(Xd_0__inst_mult_17_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_50 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[128]),
	.datac(!din_a[128]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_158 ),
	.cout(Xd_0__inst_mult_16_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_50 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[120]),
	.datac(!din_a[120]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_158 ),
	.cout(Xd_0__inst_mult_15_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_50 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[112]),
	.datac(!din_a[112]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_158 ),
	.cout(Xd_0__inst_mult_14_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_50 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[104]),
	.datac(!din_a[104]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_158 ),
	.cout(Xd_0__inst_mult_13_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_50 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[96]),
	.datac(!din_a[96]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_158 ),
	.cout(Xd_0__inst_mult_12_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_50 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[88]),
	.datac(!din_a[88]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_158 ),
	.cout(Xd_0__inst_mult_11_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_50 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[80]),
	.datac(!din_a[80]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_144 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_158 ),
	.cout(Xd_0__inst_mult_10_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_50 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[72]),
	.datac(!din_a[72]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_158 ),
	.cout(Xd_0__inst_mult_9_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_50 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[64]),
	.datac(!din_a[64]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_158 ),
	.cout(Xd_0__inst_mult_8_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_50 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[56]),
	.datac(!din_a[56]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_158 ),
	.cout(Xd_0__inst_mult_7_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_50 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[48]),
	.datac(!din_a[48]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_158 ),
	.cout(Xd_0__inst_mult_6_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_50 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[40]),
	.datac(!din_a[40]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_149 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_158 ),
	.cout(Xd_0__inst_mult_5_159 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_48 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[32]),
	.datac(!din_a[32]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_149 ),
	.cout(Xd_0__inst_mult_4_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_48 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[24]),
	.datac(!din_a[24]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_149 ),
	.cout(Xd_0__inst_mult_3_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_48 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[16]),
	.datac(!din_a[16]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_149 ),
	.cout(Xd_0__inst_mult_2_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_48 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[8]),
	.datac(!din_a[8]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_149 ),
	.cout(Xd_0__inst_mult_1_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_48 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[0]),
	.datac(!din_a[0]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_140 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_149 ),
	.cout(Xd_0__inst_mult_0_150 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_154 ),
	.cout(Xd_0__inst_mult_23_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_154 ),
	.cout(Xd_0__inst_mult_22_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_154 ),
	.cout(Xd_0__inst_mult_21_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_163 ),
	.cout(Xd_0__inst_mult_20_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_154 ),
	.cout(Xd_0__inst_mult_25_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_163 ),
	.cout(Xd_0__inst_mult_19_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_163 ),
	.cout(Xd_0__inst_mult_18_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_163 ),
	.cout(Xd_0__inst_mult_17_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_154 ),
	.cout(Xd_0__inst_mult_24_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_154 ),
	.cout(Xd_0__inst_mult_4_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_154 ),
	.cout(Xd_0__inst_mult_26_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_163 ),
	.cout(Xd_0__inst_mult_16_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_163 ),
	.cout(Xd_0__inst_mult_12_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_50 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_159 ),
	.cout(Xd_0__inst_mult_23_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_163 ),
	.cout(Xd_0__inst_mult_5_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_163 ),
	.cout(Xd_0__inst_mult_6_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_163 ),
	.cout(Xd_0__inst_mult_7_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_163 ),
	.cout(Xd_0__inst_mult_8_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_163 ),
	.cout(Xd_0__inst_mult_9_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_52 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_168 ),
	.cout(Xd_0__inst_mult_19_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_163 ),
	.cout(Xd_0__inst_mult_10_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_163 ),
	.cout(Xd_0__inst_mult_11_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_163 ),
	.cout(Xd_0__inst_mult_13_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_163 ),
	.cout(Xd_0__inst_mult_14_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_163 ),
	.cout(Xd_0__inst_mult_15_164 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_52 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_168 ),
	.cout(Xd_0__inst_mult_16_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_52 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_168 ),
	.cout(Xd_0__inst_mult_17_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_52 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_168 ),
	.cout(Xd_0__inst_mult_18_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_154 ),
	.cout(Xd_0__inst_mult_30_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_52 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_168 ),
	.cout(Xd_0__inst_mult_20_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_50 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_159 ),
	.cout(Xd_0__inst_mult_21_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_50 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_159 ),
	.cout(Xd_0__inst_mult_22_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_52 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[45]),
	.datac(!din_a[43]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_168 ),
	.cout(Xd_0__inst_mult_5_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_52 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[53]),
	.datac(!din_a[51]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_168 ),
	.cout(Xd_0__inst_mult_6_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_52 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[61]),
	.datac(!din_a[59]),
	.datad(!din_b[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_168 ),
	.cout(Xd_0__inst_mult_7_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_52 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[69]),
	.datac(!din_a[67]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_168 ),
	.cout(Xd_0__inst_mult_8_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_52 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[77]),
	.datac(!din_a[75]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_168 ),
	.cout(Xd_0__inst_mult_9_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_53 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[165]),
	.datac(!din_a[163]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_173 ),
	.cout(Xd_0__inst_mult_20_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_53 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[157]),
	.datac(!din_a[155]),
	.datad(!din_b[155]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_173 ),
	.cout(Xd_0__inst_mult_19_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_52 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[93]),
	.datac(!din_a[91]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_168 ),
	.cout(Xd_0__inst_mult_11_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_53 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[149]),
	.datac(!din_a[147]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_173 ),
	.cout(Xd_0__inst_mult_18_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_53 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[141]),
	.datac(!din_a[139]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_173 ),
	.cout(Xd_0__inst_mult_17_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_53 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[133]),
	.datac(!din_a[131]),
	.datad(!din_b[131]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_173 ),
	.cout(Xd_0__inst_mult_16_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_52 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[85]),
	.datac(!din_a[83]),
	.datad(!din_b[83]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_168 ),
	.cout(Xd_0__inst_mult_10_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_52 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[125]),
	.datac(!din_a[123]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_168 ),
	.cout(Xd_0__inst_mult_15_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_52 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[117]),
	.datac(!din_a[115]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_168 ),
	.cout(Xd_0__inst_mult_14_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_52 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[109]),
	.datac(!din_a[107]),
	.datad(!din_b[107]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_168 ),
	.cout(Xd_0__inst_mult_13_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_23 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_23_sumout ),
	.cout(Xd_0__inst_mult_16_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_52 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[101]),
	.datac(!din_a[99]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_168 ),
	.cout(Xd_0__inst_mult_12_169 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_53 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_173 ),
	.cout(Xd_0__inst_mult_15_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_28 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[190]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_28_sumout ),
	.cout(Xd_0__inst_mult_23_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_50 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_159 ),
	.cout(Xd_0__inst_mult_30_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_28 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[182]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_28_sumout ),
	.cout(Xd_0__inst_mult_22_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_154 ),
	.cout(Xd_0__inst_mult_28_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_23 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[5]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_23_sumout ),
	.cout(Xd_0__inst_mult_0_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_154 ),
	.cout(Xd_0__inst_mult_0_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_50 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_159 ),
	.cout(Xd_0__inst_mult_26_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_28 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_28_sumout ),
	.cout(Xd_0__inst_mult_5_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_154 ),
	.cout(Xd_0__inst_mult_3_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_28 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[133]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_28_sumout ),
	.cout(Xd_0__inst_mult_16_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_49 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_154 ),
	.cout(Xd_0__inst_mult_1_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_49 (
// Equation(s):

	.dataa(!din_a[251]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_31_239 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_154 ),
	.cout(Xd_0__inst_mult_31_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_31_50 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[251]),
	.datac(!din_a[249]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_159 ),
	.cout(Xd_0__inst_mult_31_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_51 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[189]),
	.datac(!din_a[188]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_164 ),
	.cout(Xd_0__inst_mult_23_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_51 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[240]),
	.datac(!Xd_0__inst_mult_30_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_164 ),
	.cout(Xd_0__inst_mult_30_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_30_52 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[243]),
	.datac(!din_a[241]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_169 ),
	.cout(Xd_0__inst_mult_30_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_51 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[181]),
	.datac(!din_a[180]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_164 ),
	.cout(Xd_0__inst_mult_22_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_49 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[232]),
	.datac(!Xd_0__inst_mult_29_239 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_154 ),
	.cout(Xd_0__inst_mult_29_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_29_50 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[235]),
	.datac(!din_a[233]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_159 ),
	.cout(Xd_0__inst_mult_29_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_51 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[173]),
	.datac(!din_a[172]),
	.datad(!din_b[174]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_164 ),
	.cout(Xd_0__inst_mult_21_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_50 (
// Equation(s):

	.dataa(!din_a[227]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_28_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_159 ),
	.cout(Xd_0__inst_mult_28_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_28_51 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[227]),
	.datac(!din_a[225]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_164 ),
	.cout(Xd_0__inst_mult_28_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_54 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[165]),
	.datac(!din_a[164]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_178 ),
	.cout(Xd_0__inst_mult_20_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_49 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[216]),
	.datac(!Xd_0__inst_mult_27_239 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_154 ),
	.cout(Xd_0__inst_mult_27_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_27_50 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[219]),
	.datac(!din_a[217]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_159 ),
	.cout(Xd_0__inst_mult_27_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_50 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[205]),
	.datac(!din_a[204]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_159 ),
	.cout(Xd_0__inst_mult_25_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_51 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[208]),
	.datac(!Xd_0__inst_mult_26_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_164 ),
	.cout(Xd_0__inst_mult_26_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_26_52 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[211]),
	.datac(!din_a[209]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_169 ),
	.cout(Xd_0__inst_mult_26_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_54 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[157]),
	.datac(!din_a[156]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_178 ),
	.cout(Xd_0__inst_mult_19_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_51 (
// Equation(s):

	.dataa(!din_a[203]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_25_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_164 ),
	.cout(Xd_0__inst_mult_25_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_25_52 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[203]),
	.datac(!din_a[201]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_169 ),
	.cout(Xd_0__inst_mult_25_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_54 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[149]),
	.datac(!din_a[148]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_178 ),
	.cout(Xd_0__inst_mult_18_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_50 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[192]),
	.datac(!Xd_0__inst_mult_24_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_159 ),
	.cout(Xd_0__inst_mult_24_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_24_51 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[195]),
	.datac(!din_a[193]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_164 ),
	.cout(Xd_0__inst_mult_24_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_54 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[141]),
	.datac(!din_a[140]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_178 ),
	.cout(Xd_0__inst_mult_17_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_52 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[184]),
	.datac(!Xd_0__inst_mult_23_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_169 ),
	.cout(Xd_0__inst_mult_23_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_23_53 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[187]),
	.datac(!din_a[185]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_174 ),
	.cout(Xd_0__inst_mult_23_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_52 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[197]),
	.datac(!din_a[196]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_169 ),
	.cout(Xd_0__inst_mult_24_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_52 (
// Equation(s):

	.dataa(!din_a[179]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_22_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_169 ),
	.cout(Xd_0__inst_mult_22_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_22_53 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[179]),
	.datac(!din_a[177]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_174 ),
	.cout(Xd_0__inst_mult_22_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_50 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_159 ),
	.cout(Xd_0__inst_mult_4_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_52 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[168]),
	.datac(!Xd_0__inst_mult_21_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_169 ),
	.cout(Xd_0__inst_mult_21_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_21_53 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[171]),
	.datac(!din_a[169]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_174 ),
	.cout(Xd_0__inst_mult_21_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_53 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[213]),
	.datac(!din_a[212]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_174 ),
	.cout(Xd_0__inst_mult_26_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_55 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[160]),
	.datac(!Xd_0__inst_mult_20_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_183 ),
	.cout(Xd_0__inst_mult_20_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_20_56 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[163]),
	.datac(!din_a[161]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_188 ),
	.cout(Xd_0__inst_mult_20_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_54 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[133]),
	.datac(!din_a[132]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_178 ),
	.cout(Xd_0__inst_mult_16_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_55 (
// Equation(s):

	.dataa(!din_a[155]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_19_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_183 ),
	.cout(Xd_0__inst_mult_19_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_19_56 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[155]),
	.datac(!din_a[153]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_188 ),
	.cout(Xd_0__inst_mult_19_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_53 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[98]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_173 ),
	.cout(Xd_0__inst_mult_12_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_55 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[144]),
	.datac(!Xd_0__inst_mult_18_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_183 ),
	.cout(Xd_0__inst_mult_18_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_18_56 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[147]),
	.datac(!din_a[145]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_188 ),
	.cout(Xd_0__inst_mult_18_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_54 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[186]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_179 ),
	.cout(Xd_0__inst_mult_23_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_55 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[136]),
	.datac(!Xd_0__inst_mult_17_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_183 ),
	.cout(Xd_0__inst_mult_17_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_17_56 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[139]),
	.datac(!din_a[137]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_188 ),
	.cout(Xd_0__inst_mult_17_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_53 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[42]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_173 ),
	.cout(Xd_0__inst_mult_5_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_55 (
// Equation(s):

	.dataa(!din_a[131]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_16_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_183 ),
	.cout(Xd_0__inst_mult_16_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_16_56 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[131]),
	.datac(!din_a[129]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_188 ),
	.cout(Xd_0__inst_mult_16_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_53 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[50]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_173 ),
	.cout(Xd_0__inst_mult_6_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_54 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[120]),
	.datac(!Xd_0__inst_mult_15_273 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_178 ),
	.cout(Xd_0__inst_mult_15_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_15_55 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[123]),
	.datac(!din_a[121]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_183 ),
	.cout(Xd_0__inst_mult_15_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_53 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_173 ),
	.cout(Xd_0__inst_mult_7_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_53 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[112]),
	.datac(!Xd_0__inst_mult_14_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_173 ),
	.cout(Xd_0__inst_mult_14_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_14_54 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[115]),
	.datac(!din_a[113]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_178 ),
	.cout(Xd_0__inst_mult_14_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_53 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[66]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_173 ),
	.cout(Xd_0__inst_mult_8_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_53 (
// Equation(s):

	.dataa(!din_a[107]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_13_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_173 ),
	.cout(Xd_0__inst_mult_13_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_13_54 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[107]),
	.datac(!din_a[105]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_178 ),
	.cout(Xd_0__inst_mult_13_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_53 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[74]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_173 ),
	.cout(Xd_0__inst_mult_9_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_54 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[96]),
	.datac(!Xd_0__inst_mult_12_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_178 ),
	.cout(Xd_0__inst_mult_12_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_12_55 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[99]),
	.datac(!din_a[97]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_183 ),
	.cout(Xd_0__inst_mult_12_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_57 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[154]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_193 ),
	.cout(Xd_0__inst_mult_19_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_53 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[88]),
	.datac(!Xd_0__inst_mult_11_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_173 ),
	.cout(Xd_0__inst_mult_11_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_11_54 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[91]),
	.datac(!din_a[89]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_178 ),
	.cout(Xd_0__inst_mult_11_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_53 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_173 ),
	.cout(Xd_0__inst_mult_10_174 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_54 (
// Equation(s):

	.dataa(!din_a[83]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_10_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_178 ),
	.cout(Xd_0__inst_mult_10_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_10_55 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[83]),
	.datac(!din_a[81]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_183 ),
	.cout(Xd_0__inst_mult_10_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_55 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_183 ),
	.cout(Xd_0__inst_mult_11_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_54 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[72]),
	.datac(!Xd_0__inst_mult_9_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_178 ),
	.cout(Xd_0__inst_mult_9_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_9_55 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[75]),
	.datac(!din_a[73]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_183 ),
	.cout(Xd_0__inst_mult_9_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_55 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[106]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_183 ),
	.cout(Xd_0__inst_mult_13_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_54 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[64]),
	.datac(!Xd_0__inst_mult_8_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_178 ),
	.cout(Xd_0__inst_mult_8_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_8_55 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[67]),
	.datac(!din_a[65]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_183 ),
	.cout(Xd_0__inst_mult_8_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_55 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[114]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_183 ),
	.cout(Xd_0__inst_mult_14_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_54 (
// Equation(s):

	.dataa(!din_a[59]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_7_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_178 ),
	.cout(Xd_0__inst_mult_7_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_7_55 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[59]),
	.datac(!din_a[57]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_183 ),
	.cout(Xd_0__inst_mult_7_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_56 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[122]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_188 ),
	.cout(Xd_0__inst_mult_15_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_54 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[48]),
	.datac(!Xd_0__inst_mult_6_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_178 ),
	.cout(Xd_0__inst_mult_6_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_6_55 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[51]),
	.datac(!din_a[49]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_183 ),
	.cout(Xd_0__inst_mult_6_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_57 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_193 ),
	.cout(Xd_0__inst_mult_16_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_54 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[40]),
	.datac(!Xd_0__inst_mult_5_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_178 ),
	.cout(Xd_0__inst_mult_5_179 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_5_55 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[43]),
	.datac(!din_a[41]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_183 ),
	.cout(Xd_0__inst_mult_5_184 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_57 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[138]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_193 ),
	.cout(Xd_0__inst_mult_17_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_51 (
// Equation(s):

	.dataa(!din_a[35]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_4_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_164 ),
	.cout(Xd_0__inst_mult_4_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_4_52 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[35]),
	.datac(!din_a[33]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_169 ),
	.cout(Xd_0__inst_mult_4_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_57 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[146]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_193 ),
	.cout(Xd_0__inst_mult_18_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_50 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[24]),
	.datac(!Xd_0__inst_mult_3_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_159 ),
	.cout(Xd_0__inst_mult_3_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_3_51 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[27]),
	.datac(!din_a[25]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_164 ),
	.cout(Xd_0__inst_mult_3_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_53 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[245]),
	.datac(!din_a[244]),
	.datad(!din_b[246]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_174 ),
	.cout(Xd_0__inst_mult_30_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_49 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[16]),
	.datac(!Xd_0__inst_mult_2_239 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_154 ),
	.cout(Xd_0__inst_mult_2_155 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_2_50 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[19]),
	.datac(!din_a[17]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_159 ),
	.cout(Xd_0__inst_mult_2_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_57 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[162]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_193 ),
	.cout(Xd_0__inst_mult_20_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_50 (
// Equation(s):

	.dataa(!din_a[11]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_1_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_159 ),
	.cout(Xd_0__inst_mult_1_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_1_51 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[11]),
	.datac(!din_a[9]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_164 ),
	.cout(Xd_0__inst_mult_1_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_54 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[170]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_179 ),
	.cout(Xd_0__inst_mult_21_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_50 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[0]),
	.datac(!Xd_0__inst_mult_0_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_159 ),
	.cout(Xd_0__inst_mult_0_160 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_0_51 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[3]),
	.datac(!din_a[1]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_164 ),
	.cout(Xd_0__inst_mult_0_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_54 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[178]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_179 ),
	.cout(Xd_0__inst_mult_22_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_51 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_31_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_164 ),
	.cout(Xd_0__inst_mult_31_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_52 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[251]),
	.datac(!din_a[248]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_169 ),
	.cout(Xd_0__inst_mult_31_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_54 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[240]),
	.datac(!Xd_0__inst_mult_30_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_179 ),
	.cout(Xd_0__inst_mult_30_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_55 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[243]),
	.datac(!din_a[240]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_184 ),
	.cout(Xd_0__inst_mult_30_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_51 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[232]),
	.datac(!Xd_0__inst_mult_29_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_164 ),
	.cout(Xd_0__inst_mult_29_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_52 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[235]),
	.datac(!din_a[232]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_169 ),
	.cout(Xd_0__inst_mult_29_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_52 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_28_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_169 ),
	.cout(Xd_0__inst_mult_28_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_53 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[227]),
	.datac(!din_a[224]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_174 ),
	.cout(Xd_0__inst_mult_28_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_51 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[216]),
	.datac(!Xd_0__inst_mult_27_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_164 ),
	.cout(Xd_0__inst_mult_27_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_52 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[219]),
	.datac(!din_a[216]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_169 ),
	.cout(Xd_0__inst_mult_27_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_54 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[208]),
	.datac(!Xd_0__inst_mult_26_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_179 ),
	.cout(Xd_0__inst_mult_26_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_55 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[211]),
	.datac(!din_a[208]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_184 ),
	.cout(Xd_0__inst_mult_26_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_53 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_25_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_174 ),
	.cout(Xd_0__inst_mult_25_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_54 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[203]),
	.datac(!din_a[200]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_179 ),
	.cout(Xd_0__inst_mult_25_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_53 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[192]),
	.datac(!Xd_0__inst_mult_24_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_174 ),
	.cout(Xd_0__inst_mult_24_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_54 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[195]),
	.datac(!din_a[192]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_179 ),
	.cout(Xd_0__inst_mult_24_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_55 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[184]),
	.datac(!Xd_0__inst_mult_23_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_184 ),
	.cout(Xd_0__inst_mult_23_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_56 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[187]),
	.datac(!din_a[184]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_189 ),
	.cout(Xd_0__inst_mult_23_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_55 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_22_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_184 ),
	.cout(Xd_0__inst_mult_22_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_56 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[179]),
	.datac(!din_a[176]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_189 ),
	.cout(Xd_0__inst_mult_22_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_55 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[168]),
	.datac(!Xd_0__inst_mult_21_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_184 ),
	.cout(Xd_0__inst_mult_21_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_56 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[171]),
	.datac(!din_a[168]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_189 ),
	.cout(Xd_0__inst_mult_21_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_58 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[160]),
	.datac(!Xd_0__inst_mult_20_293 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_198 ),
	.cout(Xd_0__inst_mult_20_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_59 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[163]),
	.datac(!din_a[160]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_203 ),
	.cout(Xd_0__inst_mult_20_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_58 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_19_293 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_198 ),
	.cout(Xd_0__inst_mult_19_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_59 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[155]),
	.datac(!din_a[152]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_203 ),
	.cout(Xd_0__inst_mult_19_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_58 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[144]),
	.datac(!Xd_0__inst_mult_18_293 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_198 ),
	.cout(Xd_0__inst_mult_18_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_59 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[147]),
	.datac(!din_a[144]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_203 ),
	.cout(Xd_0__inst_mult_18_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_58 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[136]),
	.datac(!Xd_0__inst_mult_17_293 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_198 ),
	.cout(Xd_0__inst_mult_17_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_59 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[139]),
	.datac(!din_a[136]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_203 ),
	.cout(Xd_0__inst_mult_17_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_58 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_16_293 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_198 ),
	.cout(Xd_0__inst_mult_16_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_59 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[131]),
	.datac(!din_a[128]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_203 ),
	.cout(Xd_0__inst_mult_16_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_57 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[120]),
	.datac(!Xd_0__inst_mult_15_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_193 ),
	.cout(Xd_0__inst_mult_15_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_58 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[123]),
	.datac(!din_a[120]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_198 ),
	.cout(Xd_0__inst_mult_15_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_56 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[112]),
	.datac(!Xd_0__inst_mult_14_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_188 ),
	.cout(Xd_0__inst_mult_14_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_57 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[115]),
	.datac(!din_a[112]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_193 ),
	.cout(Xd_0__inst_mult_14_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_56 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_13_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_188 ),
	.cout(Xd_0__inst_mult_13_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_57 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[107]),
	.datac(!din_a[104]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_193 ),
	.cout(Xd_0__inst_mult_13_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_56 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[96]),
	.datac(!Xd_0__inst_mult_12_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_188 ),
	.cout(Xd_0__inst_mult_12_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_57 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[99]),
	.datac(!din_a[96]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_193 ),
	.cout(Xd_0__inst_mult_12_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_56 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[88]),
	.datac(!Xd_0__inst_mult_11_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_174 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_188 ),
	.cout(Xd_0__inst_mult_11_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_57 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[91]),
	.datac(!din_a[88]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_193 ),
	.cout(Xd_0__inst_mult_11_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_56 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_10_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_188 ),
	.cout(Xd_0__inst_mult_10_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_57 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[83]),
	.datac(!din_a[80]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_193 ),
	.cout(Xd_0__inst_mult_10_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_56 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[72]),
	.datac(!Xd_0__inst_mult_9_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_188 ),
	.cout(Xd_0__inst_mult_9_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_57 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[75]),
	.datac(!din_a[72]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_193 ),
	.cout(Xd_0__inst_mult_9_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_56 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[64]),
	.datac(!Xd_0__inst_mult_8_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_188 ),
	.cout(Xd_0__inst_mult_8_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_57 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[67]),
	.datac(!din_a[64]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_193 ),
	.cout(Xd_0__inst_mult_8_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_56 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_7_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_188 ),
	.cout(Xd_0__inst_mult_7_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_57 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[59]),
	.datac(!din_a[56]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_193 ),
	.cout(Xd_0__inst_mult_7_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_56 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[48]),
	.datac(!Xd_0__inst_mult_6_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_188 ),
	.cout(Xd_0__inst_mult_6_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_57 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[51]),
	.datac(!din_a[48]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_193 ),
	.cout(Xd_0__inst_mult_6_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_56 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[40]),
	.datac(!Xd_0__inst_mult_5_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_188 ),
	.cout(Xd_0__inst_mult_5_189 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_57 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[43]),
	.datac(!din_a[40]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_193 ),
	.cout(Xd_0__inst_mult_5_194 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_53 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_4_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_174 ),
	.cout(Xd_0__inst_mult_4_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_54 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[35]),
	.datac(!din_a[32]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_179 ),
	.cout(Xd_0__inst_mult_4_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_52 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[24]),
	.datac(!Xd_0__inst_mult_3_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_169 ),
	.cout(Xd_0__inst_mult_3_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_53 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[27]),
	.datac(!din_a[24]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_174 ),
	.cout(Xd_0__inst_mult_3_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_51 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[16]),
	.datac(!Xd_0__inst_mult_2_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_155 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_164 ),
	.cout(Xd_0__inst_mult_2_165 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_52 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[19]),
	.datac(!din_a[16]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_169 ),
	.cout(Xd_0__inst_mult_2_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_52 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_1_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_169 ),
	.cout(Xd_0__inst_mult_1_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_53 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[11]),
	.datac(!din_a[8]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_174 ),
	.cout(Xd_0__inst_mult_1_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_52 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[0]),
	.datac(!Xd_0__inst_mult_0_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_169 ),
	.cout(Xd_0__inst_mult_0_170 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_53 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[3]),
	.datac(!din_a[0]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_174 ),
	.cout(Xd_0__inst_mult_0_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_53 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_31_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_174 ),
	.cout(Xd_0__inst_mult_31_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_54 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[251]),
	.datac(!din_a[248]),
	.datad(!din_b[253]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_179 ),
	.cout(Xd_0__inst_mult_31_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_56 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[240]),
	.datac(!Xd_0__inst_mult_30_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_189 ),
	.cout(Xd_0__inst_mult_30_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_57 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[243]),
	.datac(!din_a[240]),
	.datad(!din_b[245]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_194 ),
	.cout(Xd_0__inst_mult_30_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_53 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[232]),
	.datac(!Xd_0__inst_mult_29_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_174 ),
	.cout(Xd_0__inst_mult_29_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_54 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[235]),
	.datac(!din_a[232]),
	.datad(!din_b[237]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_179 ),
	.cout(Xd_0__inst_mult_29_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_54 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_28_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_179 ),
	.cout(Xd_0__inst_mult_28_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_55 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[227]),
	.datac(!din_a[224]),
	.datad(!din_b[229]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_184 ),
	.cout(Xd_0__inst_mult_28_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_53 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[216]),
	.datac(!Xd_0__inst_mult_27_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_174 ),
	.cout(Xd_0__inst_mult_27_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_54 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[219]),
	.datac(!din_a[216]),
	.datad(!din_b[221]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_179 ),
	.cout(Xd_0__inst_mult_27_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_56 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[208]),
	.datac(!Xd_0__inst_mult_26_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_189 ),
	.cout(Xd_0__inst_mult_26_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_57 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[211]),
	.datac(!din_a[208]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_194 ),
	.cout(Xd_0__inst_mult_26_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_55 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_25_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_184 ),
	.cout(Xd_0__inst_mult_25_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_56 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[203]),
	.datac(!din_a[200]),
	.datad(!din_b[205]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_189 ),
	.cout(Xd_0__inst_mult_25_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_55 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[192]),
	.datac(!Xd_0__inst_mult_24_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_184 ),
	.cout(Xd_0__inst_mult_24_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_56 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[195]),
	.datac(!din_a[192]),
	.datad(!din_b[197]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_189 ),
	.cout(Xd_0__inst_mult_24_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_57 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[184]),
	.datac(!Xd_0__inst_mult_23_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_194 ),
	.cout(Xd_0__inst_mult_23_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_58 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[187]),
	.datac(!din_a[184]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_199 ),
	.cout(Xd_0__inst_mult_23_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_57 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_22_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_194 ),
	.cout(Xd_0__inst_mult_22_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_58 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[179]),
	.datac(!din_a[176]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_199 ),
	.cout(Xd_0__inst_mult_22_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_57 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[168]),
	.datac(!Xd_0__inst_mult_21_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_194 ),
	.cout(Xd_0__inst_mult_21_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_58 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[171]),
	.datac(!din_a[168]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_199 ),
	.cout(Xd_0__inst_mult_21_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_60 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[160]),
	.datac(!Xd_0__inst_mult_20_298 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_208 ),
	.cout(Xd_0__inst_mult_20_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_61 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[163]),
	.datac(!din_a[160]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_213 ),
	.cout(Xd_0__inst_mult_20_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_60 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_19_298 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_208 ),
	.cout(Xd_0__inst_mult_19_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_61 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[155]),
	.datac(!din_a[152]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_213 ),
	.cout(Xd_0__inst_mult_19_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_60 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[144]),
	.datac(!Xd_0__inst_mult_18_298 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_208 ),
	.cout(Xd_0__inst_mult_18_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_61 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[147]),
	.datac(!din_a[144]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_213 ),
	.cout(Xd_0__inst_mult_18_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_60 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[136]),
	.datac(!Xd_0__inst_mult_17_298 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_208 ),
	.cout(Xd_0__inst_mult_17_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_61 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[139]),
	.datac(!din_a[136]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_213 ),
	.cout(Xd_0__inst_mult_17_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_60 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_16_298 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_208 ),
	.cout(Xd_0__inst_mult_16_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_61 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[131]),
	.datac(!din_a[128]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_213 ),
	.cout(Xd_0__inst_mult_16_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_59 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[120]),
	.datac(!Xd_0__inst_mult_15_293 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_194 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_203 ),
	.cout(Xd_0__inst_mult_15_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_60 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[123]),
	.datac(!din_a[120]),
	.datad(!din_b[125]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_208 ),
	.cout(Xd_0__inst_mult_15_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_58 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[112]),
	.datac(!Xd_0__inst_mult_14_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_198 ),
	.cout(Xd_0__inst_mult_14_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_59 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[115]),
	.datac(!din_a[112]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_203 ),
	.cout(Xd_0__inst_mult_14_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_58 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_13_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_198 ),
	.cout(Xd_0__inst_mult_13_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_59 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[107]),
	.datac(!din_a[104]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_203 ),
	.cout(Xd_0__inst_mult_13_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_58 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[96]),
	.datac(!Xd_0__inst_mult_12_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_198 ),
	.cout(Xd_0__inst_mult_12_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_59 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[99]),
	.datac(!din_a[96]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_203 ),
	.cout(Xd_0__inst_mult_12_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_58 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[88]),
	.datac(!Xd_0__inst_mult_11_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_198 ),
	.cout(Xd_0__inst_mult_11_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_59 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[91]),
	.datac(!din_a[88]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_179 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_203 ),
	.cout(Xd_0__inst_mult_11_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_58 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_10_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_198 ),
	.cout(Xd_0__inst_mult_10_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_59 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[83]),
	.datac(!din_a[80]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_203 ),
	.cout(Xd_0__inst_mult_10_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_58 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[72]),
	.datac(!Xd_0__inst_mult_9_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_198 ),
	.cout(Xd_0__inst_mult_9_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_59 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[75]),
	.datac(!din_a[72]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_203 ),
	.cout(Xd_0__inst_mult_9_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_58 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[64]),
	.datac(!Xd_0__inst_mult_8_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_198 ),
	.cout(Xd_0__inst_mult_8_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_59 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[67]),
	.datac(!din_a[64]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_203 ),
	.cout(Xd_0__inst_mult_8_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_58 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_7_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_198 ),
	.cout(Xd_0__inst_mult_7_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_59 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[59]),
	.datac(!din_a[56]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_203 ),
	.cout(Xd_0__inst_mult_7_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_58 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[48]),
	.datac(!Xd_0__inst_mult_6_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_198 ),
	.cout(Xd_0__inst_mult_6_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_59 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[51]),
	.datac(!din_a[48]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_203 ),
	.cout(Xd_0__inst_mult_6_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_58 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[40]),
	.datac(!Xd_0__inst_mult_5_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_189 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_198 ),
	.cout(Xd_0__inst_mult_5_199 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_59 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[43]),
	.datac(!din_a[40]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_184 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_203 ),
	.cout(Xd_0__inst_mult_5_204 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_55 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_4_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_184 ),
	.cout(Xd_0__inst_mult_4_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_56 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[35]),
	.datac(!din_a[32]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_189 ),
	.cout(Xd_0__inst_mult_4_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_54 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[24]),
	.datac(!Xd_0__inst_mult_3_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_179 ),
	.cout(Xd_0__inst_mult_3_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_55 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[27]),
	.datac(!din_a[24]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_184 ),
	.cout(Xd_0__inst_mult_3_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_53 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[16]),
	.datac(!Xd_0__inst_mult_2_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_174 ),
	.cout(Xd_0__inst_mult_2_175 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_54 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[19]),
	.datac(!din_a[16]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_160 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_179 ),
	.cout(Xd_0__inst_mult_2_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_54 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_1_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_179 ),
	.cout(Xd_0__inst_mult_1_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_55 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[11]),
	.datac(!din_a[8]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_184 ),
	.cout(Xd_0__inst_mult_1_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_54 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[0]),
	.datac(!Xd_0__inst_mult_0_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_170 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_179 ),
	.cout(Xd_0__inst_mult_0_180 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_55 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[3]),
	.datac(!din_a[0]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_165 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_184 ),
	.cout(Xd_0__inst_mult_0_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_55 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_31_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_184 ),
	.cout(Xd_0__inst_mult_31_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_56 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_269 ),
	.datab(!Xd_0__inst_mult_31_274 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_189 ),
	.cout(Xd_0__inst_mult_31_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_58 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[240]),
	.datac(!Xd_0__inst_mult_30_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_199 ),
	.cout(Xd_0__inst_mult_30_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_59 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_289 ),
	.datab(!Xd_0__inst_mult_30_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_204 ),
	.cout(Xd_0__inst_mult_30_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_55 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[232]),
	.datac(!Xd_0__inst_mult_29_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_184 ),
	.cout(Xd_0__inst_mult_29_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_56 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_264 ),
	.datab(!Xd_0__inst_mult_29_269 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_189 ),
	.cout(Xd_0__inst_mult_29_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_56 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_28_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_189 ),
	.cout(Xd_0__inst_mult_28_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_57 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_279 ),
	.datab(!Xd_0__inst_mult_28_284 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_194 ),
	.cout(Xd_0__inst_mult_28_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_55 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[216]),
	.datac(!Xd_0__inst_mult_27_259 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_184 ),
	.cout(Xd_0__inst_mult_27_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_56 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_264 ),
	.datab(!Xd_0__inst_mult_27_269 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_189 ),
	.cout(Xd_0__inst_mult_27_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_58 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[208]),
	.datac(!Xd_0__inst_mult_26_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_199 ),
	.cout(Xd_0__inst_mult_26_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_59 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_289 ),
	.datab(!Xd_0__inst_mult_26_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_204 ),
	.cout(Xd_0__inst_mult_26_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_57 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_25_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_194 ),
	.cout(Xd_0__inst_mult_25_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_279 ),
	.datab(!Xd_0__inst_mult_25_284 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_199 ),
	.cout(Xd_0__inst_mult_25_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_57 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[192]),
	.datac(!Xd_0__inst_mult_24_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_194 ),
	.cout(Xd_0__inst_mult_24_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_279 ),
	.datab(!Xd_0__inst_mult_24_284 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_199 ),
	.cout(Xd_0__inst_mult_24_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_59 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[184]),
	.datac(!Xd_0__inst_mult_23_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_204 ),
	.cout(Xd_0__inst_mult_23_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_289 ),
	.datab(!Xd_0__inst_mult_23_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_209 ),
	.cout(Xd_0__inst_mult_23_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_59 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_22_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_204 ),
	.cout(Xd_0__inst_mult_22_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_289 ),
	.datab(!Xd_0__inst_mult_22_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_209 ),
	.cout(Xd_0__inst_mult_22_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_59 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[168]),
	.datac(!Xd_0__inst_mult_21_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_204 ),
	.cout(Xd_0__inst_mult_21_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_289 ),
	.datab(!Xd_0__inst_mult_21_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_209 ),
	.cout(Xd_0__inst_mult_21_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_62 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[160]),
	.datac(!Xd_0__inst_mult_20_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_218 ),
	.cout(Xd_0__inst_mult_20_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_303 ),
	.datab(!Xd_0__inst_mult_20_173 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_223 ),
	.cout(Xd_0__inst_mult_20_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_62 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_19_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_218 ),
	.cout(Xd_0__inst_mult_19_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_303 ),
	.datab(!Xd_0__inst_mult_19_173 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_223 ),
	.cout(Xd_0__inst_mult_19_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_62 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[144]),
	.datac(!Xd_0__inst_mult_18_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_218 ),
	.cout(Xd_0__inst_mult_18_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_303 ),
	.datab(!Xd_0__inst_mult_18_173 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_223 ),
	.cout(Xd_0__inst_mult_18_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_62 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[136]),
	.datac(!Xd_0__inst_mult_17_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_218 ),
	.cout(Xd_0__inst_mult_17_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_303 ),
	.datab(!Xd_0__inst_mult_17_173 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_223 ),
	.cout(Xd_0__inst_mult_17_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_62 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_16_288 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_218 ),
	.cout(Xd_0__inst_mult_16_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_303 ),
	.datab(!Xd_0__inst_mult_16_173 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_223 ),
	.cout(Xd_0__inst_mult_16_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_61 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[120]),
	.datac(!Xd_0__inst_mult_15_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_213 ),
	.cout(Xd_0__inst_mult_15_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_298 ),
	.datab(!Xd_0__inst_mult_15_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_218 ),
	.cout(Xd_0__inst_mult_15_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_60 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[112]),
	.datac(!Xd_0__inst_mult_14_273 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_208 ),
	.cout(Xd_0__inst_mult_14_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_288 ),
	.datab(!Xd_0__inst_mult_14_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_213 ),
	.cout(Xd_0__inst_mult_14_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_60 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_13_273 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_208 ),
	.cout(Xd_0__inst_mult_13_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_293 ),
	.datab(!Xd_0__inst_mult_13_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_213 ),
	.cout(Xd_0__inst_mult_13_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_60 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[96]),
	.datac(!Xd_0__inst_mult_12_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_208 ),
	.cout(Xd_0__inst_mult_12_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_288 ),
	.datab(!Xd_0__inst_mult_12_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_213 ),
	.cout(Xd_0__inst_mult_12_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_60 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[88]),
	.datac(!Xd_0__inst_mult_11_273 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_208 ),
	.cout(Xd_0__inst_mult_11_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_293 ),
	.datab(!Xd_0__inst_mult_11_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_213 ),
	.cout(Xd_0__inst_mult_11_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_60 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_10_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_208 ),
	.cout(Xd_0__inst_mult_10_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_293 ),
	.datab(!Xd_0__inst_mult_10_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_213 ),
	.cout(Xd_0__inst_mult_10_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_60 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[72]),
	.datac(!Xd_0__inst_mult_9_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_208 ),
	.cout(Xd_0__inst_mult_9_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_288 ),
	.datab(!Xd_0__inst_mult_9_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_213 ),
	.cout(Xd_0__inst_mult_9_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_60 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[64]),
	.datac(!Xd_0__inst_mult_8_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_208 ),
	.cout(Xd_0__inst_mult_8_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_293 ),
	.datab(!Xd_0__inst_mult_8_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_213 ),
	.cout(Xd_0__inst_mult_8_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_60 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_7_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_208 ),
	.cout(Xd_0__inst_mult_7_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_288 ),
	.datab(!Xd_0__inst_mult_7_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_213 ),
	.cout(Xd_0__inst_mult_7_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_60 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[48]),
	.datac(!Xd_0__inst_mult_6_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_208 ),
	.cout(Xd_0__inst_mult_6_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_293 ),
	.datab(!Xd_0__inst_mult_6_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_213 ),
	.cout(Xd_0__inst_mult_6_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_60 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[40]),
	.datac(!Xd_0__inst_mult_5_263 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_199 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_208 ),
	.cout(Xd_0__inst_mult_5_209 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_288 ),
	.datab(!Xd_0__inst_mult_5_168 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_213 ),
	.cout(Xd_0__inst_mult_5_214 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_57 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_4_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_194 ),
	.cout(Xd_0__inst_mult_4_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_279 ),
	.datab(!Xd_0__inst_mult_4_284 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_199 ),
	.cout(Xd_0__inst_mult_4_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_56 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[24]),
	.datac(!Xd_0__inst_mult_3_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_189 ),
	.cout(Xd_0__inst_mult_3_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_57 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_274 ),
	.datab(!Xd_0__inst_mult_3_279 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_194 ),
	.cout(Xd_0__inst_mult_3_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_55 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[16]),
	.datac(!Xd_0__inst_mult_2_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_175 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_184 ),
	.cout(Xd_0__inst_mult_2_185 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_56 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_269 ),
	.datab(!Xd_0__inst_mult_2_274 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_189 ),
	.cout(Xd_0__inst_mult_2_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_56 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_1_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_189 ),
	.cout(Xd_0__inst_mult_1_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_57 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_274 ),
	.datab(!Xd_0__inst_mult_1_279 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_194 ),
	.cout(Xd_0__inst_mult_1_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_56 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[0]),
	.datac(!Xd_0__inst_mult_0_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_189 ),
	.cout(Xd_0__inst_mult_0_190 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_57 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_274 ),
	.datab(!Xd_0__inst_mult_0_279 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_194 ),
	.cout(Xd_0__inst_mult_0_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_57 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[249]),
	.datac(!Xd_0__inst_mult_31_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_194 ),
	.cout(Xd_0__inst_mult_31_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_289 ),
	.datab(!Xd_0__inst_mult_31_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_199 ),
	.cout(Xd_0__inst_mult_31_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_60 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[241]),
	.datac(!Xd_0__inst_mult_30_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_209 ),
	.cout(Xd_0__inst_mult_30_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_304 ),
	.datab(!Xd_0__inst_mult_30_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_214 ),
	.cout(Xd_0__inst_mult_30_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_57 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_29_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_194 ),
	.cout(Xd_0__inst_mult_29_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_284 ),
	.datab(!Xd_0__inst_mult_29_289 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_199 ),
	.cout(Xd_0__inst_mult_29_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_58 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[225]),
	.datac(!Xd_0__inst_mult_28_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_199 ),
	.cout(Xd_0__inst_mult_28_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_59 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_294 ),
	.datab(!Xd_0__inst_mult_28_299 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_204 ),
	.cout(Xd_0__inst_mult_28_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_57 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[217]),
	.datac(!Xd_0__inst_mult_27_279 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_194 ),
	.cout(Xd_0__inst_mult_27_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_284 ),
	.datab(!Xd_0__inst_mult_27_289 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_199 ),
	.cout(Xd_0__inst_mult_27_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_60 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_26_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_209 ),
	.cout(Xd_0__inst_mult_26_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_304 ),
	.datab(!Xd_0__inst_mult_26_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_214 ),
	.cout(Xd_0__inst_mult_26_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_59 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[201]),
	.datac(!Xd_0__inst_mult_25_294 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_204 ),
	.cout(Xd_0__inst_mult_25_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_299 ),
	.datab(!Xd_0__inst_mult_25_304 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_209 ),
	.cout(Xd_0__inst_mult_25_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_59 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[193]),
	.datac(!Xd_0__inst_mult_24_294 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_204 ),
	.cout(Xd_0__inst_mult_24_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_299 ),
	.datab(!Xd_0__inst_mult_24_304 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_209 ),
	.cout(Xd_0__inst_mult_24_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_61 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_23_179 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_214 ),
	.cout(Xd_0__inst_mult_23_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_304 ),
	.datab(!Xd_0__inst_mult_23_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_219 ),
	.cout(Xd_0__inst_mult_23_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_61 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[177]),
	.datac(!Xd_0__inst_mult_22_179 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_214 ),
	.cout(Xd_0__inst_mult_22_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_304 ),
	.datab(!Xd_0__inst_mult_22_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_219 ),
	.cout(Xd_0__inst_mult_22_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_61 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[169]),
	.datac(!Xd_0__inst_mult_21_179 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_214 ),
	.cout(Xd_0__inst_mult_21_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_304 ),
	.datab(!Xd_0__inst_mult_21_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_219 ),
	.cout(Xd_0__inst_mult_21_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_64 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_20_193 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_228 ),
	.cout(Xd_0__inst_mult_20_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_313 ),
	.datab(!Xd_0__inst_mult_20_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_233 ),
	.cout(Xd_0__inst_mult_20_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_64 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[153]),
	.datac(!Xd_0__inst_mult_19_193 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_228 ),
	.cout(Xd_0__inst_mult_19_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_313 ),
	.datab(!Xd_0__inst_mult_19_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_233 ),
	.cout(Xd_0__inst_mult_19_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_64 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[145]),
	.datac(!Xd_0__inst_mult_18_193 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_228 ),
	.cout(Xd_0__inst_mult_18_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_313 ),
	.datab(!Xd_0__inst_mult_18_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_233 ),
	.cout(Xd_0__inst_mult_18_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_64 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_17_193 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_228 ),
	.cout(Xd_0__inst_mult_17_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_313 ),
	.datab(!Xd_0__inst_mult_17_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_233 ),
	.cout(Xd_0__inst_mult_17_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_64 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[129]),
	.datac(!Xd_0__inst_mult_16_193 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_228 ),
	.cout(Xd_0__inst_mult_16_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_313 ),
	.datab(!Xd_0__inst_mult_16_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_233 ),
	.cout(Xd_0__inst_mult_16_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_63 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[121]),
	.datac(!Xd_0__inst_mult_15_188 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_223 ),
	.cout(Xd_0__inst_mult_15_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_308 ),
	.datab(!Xd_0__inst_mult_15_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_228 ),
	.cout(Xd_0__inst_mult_15_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_62 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_14_183 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_218 ),
	.cout(Xd_0__inst_mult_14_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_298 ),
	.datab(!Xd_0__inst_mult_14_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_223 ),
	.cout(Xd_0__inst_mult_14_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_62 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[105]),
	.datac(!Xd_0__inst_mult_13_183 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_218 ),
	.cout(Xd_0__inst_mult_13_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_303 ),
	.datab(!Xd_0__inst_mult_13_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_223 ),
	.cout(Xd_0__inst_mult_13_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_62 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[97]),
	.datac(!Xd_0__inst_mult_12_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_218 ),
	.cout(Xd_0__inst_mult_12_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_298 ),
	.datab(!Xd_0__inst_mult_12_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_223 ),
	.cout(Xd_0__inst_mult_12_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_62 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_11_183 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_218 ),
	.cout(Xd_0__inst_mult_11_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_303 ),
	.datab(!Xd_0__inst_mult_11_143 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_223 ),
	.cout(Xd_0__inst_mult_11_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_62 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[81]),
	.datac(!Xd_0__inst_mult_10_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_218 ),
	.cout(Xd_0__inst_mult_10_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_303 ),
	.datab(!Xd_0__inst_mult_10_148 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_223 ),
	.cout(Xd_0__inst_mult_10_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_62 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[73]),
	.datac(!Xd_0__inst_mult_9_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_218 ),
	.cout(Xd_0__inst_mult_9_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_298 ),
	.datab(!Xd_0__inst_mult_9_143 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_223 ),
	.cout(Xd_0__inst_mult_9_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_62 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_8_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_218 ),
	.cout(Xd_0__inst_mult_8_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_303 ),
	.datab(!Xd_0__inst_mult_8_143 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_223 ),
	.cout(Xd_0__inst_mult_8_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_62 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[57]),
	.datac(!Xd_0__inst_mult_7_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_218 ),
	.cout(Xd_0__inst_mult_7_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_298 ),
	.datab(!Xd_0__inst_mult_7_143 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_223 ),
	.cout(Xd_0__inst_mult_7_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_62 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[49]),
	.datac(!Xd_0__inst_mult_6_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_218 ),
	.cout(Xd_0__inst_mult_6_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_303 ),
	.datab(!Xd_0__inst_mult_6_143 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_223 ),
	.cout(Xd_0__inst_mult_6_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_62 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_5_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_218 ),
	.cout(Xd_0__inst_mult_5_219 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_298 ),
	.datab(!Xd_0__inst_mult_5_143 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_223 ),
	.cout(Xd_0__inst_mult_5_224 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_59 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[33]),
	.datac(!Xd_0__inst_mult_4_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_204 ),
	.cout(Xd_0__inst_mult_4_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_294 ),
	.datab(!Xd_0__inst_mult_4_299 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_209 ),
	.cout(Xd_0__inst_mult_4_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_58 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[25]),
	.datac(!Xd_0__inst_mult_3_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_199 ),
	.cout(Xd_0__inst_mult_3_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_59 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_289 ),
	.datab(!Xd_0__inst_mult_3_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_204 ),
	.cout(Xd_0__inst_mult_3_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_57 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_2_284 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_194 ),
	.cout(Xd_0__inst_mult_2_195 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_58 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_289 ),
	.datab(!Xd_0__inst_mult_2_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_199 ),
	.cout(Xd_0__inst_mult_2_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_58 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[9]),
	.datac(!Xd_0__inst_mult_1_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_199 ),
	.cout(Xd_0__inst_mult_1_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_59 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_289 ),
	.datab(!Xd_0__inst_mult_1_294 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_204 ),
	.cout(Xd_0__inst_mult_1_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_58 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[1]),
	.datac(!Xd_0__inst_mult_0_289 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_199 ),
	.cout(Xd_0__inst_mult_0_200 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_59 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_294 ),
	.datab(!Xd_0__inst_mult_0_299 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_204 ),
	.cout(Xd_0__inst_mult_0_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_59 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[250]),
	.datac(!Xd_0__inst_mult_31_299 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_204 ),
	.cout(Xd_0__inst_mult_31_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_304 ),
	.datab(!Xd_0__inst_mult_31_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_209 ),
	.cout(Xd_0__inst_mult_31_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_62 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_30_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_219 ),
	.cout(Xd_0__inst_mult_30_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_314 ),
	.datab(!Xd_0__inst_mult_30_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_224 ),
	.cout(Xd_0__inst_mult_30_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_59 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[234]),
	.datac(!Xd_0__inst_mult_29_294 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_204 ),
	.cout(Xd_0__inst_mult_29_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_299 ),
	.datab(!Xd_0__inst_mult_29_304 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_209 ),
	.cout(Xd_0__inst_mult_29_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_60 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[226]),
	.datac(!Xd_0__inst_mult_28_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_209 ),
	.cout(Xd_0__inst_mult_28_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_304 ),
	.datab(!Xd_0__inst_mult_28_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_214 ),
	.cout(Xd_0__inst_mult_28_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_59 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_27_294 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_204 ),
	.cout(Xd_0__inst_mult_27_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_299 ),
	.datab(!Xd_0__inst_mult_27_304 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_209 ),
	.cout(Xd_0__inst_mult_27_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_62 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[210]),
	.datac(!Xd_0__inst_mult_26_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_219 ),
	.cout(Xd_0__inst_mult_26_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_314 ),
	.datab(!Xd_0__inst_mult_26_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_224 ),
	.cout(Xd_0__inst_mult_26_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_61 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[202]),
	.datac(!Xd_0__inst_mult_25_309 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_214 ),
	.cout(Xd_0__inst_mult_25_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_314 ),
	.datab(!Xd_0__inst_mult_25_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_219 ),
	.cout(Xd_0__inst_mult_25_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_61 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_24_309 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_214 ),
	.cout(Xd_0__inst_mult_24_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_314 ),
	.datab(!Xd_0__inst_mult_24_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_219 ),
	.cout(Xd_0__inst_mult_24_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_63 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[186]),
	.datac(!Xd_0__inst_mult_23_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_224 ),
	.cout(Xd_0__inst_mult_23_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_314 ),
	.datab(!Xd_0__inst_mult_23_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_229 ),
	.cout(Xd_0__inst_mult_23_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_63 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[178]),
	.datac(!Xd_0__inst_mult_22_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_224 ),
	.cout(Xd_0__inst_mult_22_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_314 ),
	.datab(!Xd_0__inst_mult_22_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_229 ),
	.cout(Xd_0__inst_mult_22_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_63 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_21_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_224 ),
	.cout(Xd_0__inst_mult_21_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_314 ),
	.datab(!Xd_0__inst_mult_21_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_229 ),
	.cout(Xd_0__inst_mult_21_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_66 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[162]),
	.datac(!Xd_0__inst_mult_20_168 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_238 ),
	.cout(Xd_0__inst_mult_20_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_318 ),
	.datab(!Xd_0__inst_mult_20_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_243 ),
	.cout(Xd_0__inst_mult_20_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_66 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[154]),
	.datac(!Xd_0__inst_mult_19_168 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_238 ),
	.cout(Xd_0__inst_mult_19_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_318 ),
	.datab(!Xd_0__inst_mult_19_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_243 ),
	.cout(Xd_0__inst_mult_19_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_66 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_18_168 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_238 ),
	.cout(Xd_0__inst_mult_18_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_318 ),
	.datab(!Xd_0__inst_mult_18_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_243 ),
	.cout(Xd_0__inst_mult_18_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_66 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[138]),
	.datac(!Xd_0__inst_mult_17_168 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_238 ),
	.cout(Xd_0__inst_mult_17_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_318 ),
	.datab(!Xd_0__inst_mult_17_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_243 ),
	.cout(Xd_0__inst_mult_17_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_66 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[130]),
	.datac(!Xd_0__inst_mult_16_168 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_238 ),
	.cout(Xd_0__inst_mult_16_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_318 ),
	.datab(!Xd_0__inst_mult_16_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_243 ),
	.cout(Xd_0__inst_mult_16_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_65 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_15_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_233 ),
	.cout(Xd_0__inst_mult_15_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_66 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_313 ),
	.datab(!Xd_0__inst_mult_15_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_238 ),
	.cout(Xd_0__inst_mult_15_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_64 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[114]),
	.datac(!Xd_0__inst_mult_14_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_228 ),
	.cout(Xd_0__inst_mult_14_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_303 ),
	.datab(!Xd_0__inst_mult_14_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_233 ),
	.cout(Xd_0__inst_mult_14_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_64 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[106]),
	.datac(!Xd_0__inst_mult_13_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_228 ),
	.cout(Xd_0__inst_mult_13_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_308 ),
	.datab(!Xd_0__inst_mult_13_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_233 ),
	.cout(Xd_0__inst_mult_13_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_64 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_12_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_228 ),
	.cout(Xd_0__inst_mult_12_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_303 ),
	.datab(!Xd_0__inst_mult_12_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_233 ),
	.cout(Xd_0__inst_mult_12_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_64 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[90]),
	.datac(!Xd_0__inst_mult_11_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_228 ),
	.cout(Xd_0__inst_mult_11_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_308 ),
	.datab(!Xd_0__inst_mult_11_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_233 ),
	.cout(Xd_0__inst_mult_11_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_64 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[82]),
	.datac(!Xd_0__inst_mult_10_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_228 ),
	.cout(Xd_0__inst_mult_10_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_308 ),
	.datab(!Xd_0__inst_mult_10_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_233 ),
	.cout(Xd_0__inst_mult_10_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_64 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_9_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_228 ),
	.cout(Xd_0__inst_mult_9_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_303 ),
	.datab(!Xd_0__inst_mult_9_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_233 ),
	.cout(Xd_0__inst_mult_9_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_64 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[66]),
	.datac(!Xd_0__inst_mult_8_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_228 ),
	.cout(Xd_0__inst_mult_8_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_308 ),
	.datab(!Xd_0__inst_mult_8_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_233 ),
	.cout(Xd_0__inst_mult_8_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_64 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[58]),
	.datac(!Xd_0__inst_mult_7_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_228 ),
	.cout(Xd_0__inst_mult_7_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_303 ),
	.datab(!Xd_0__inst_mult_7_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_233 ),
	.cout(Xd_0__inst_mult_7_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_64 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_6_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_228 ),
	.cout(Xd_0__inst_mult_6_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_308 ),
	.datab(!Xd_0__inst_mult_6_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_233 ),
	.cout(Xd_0__inst_mult_6_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_64 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[42]),
	.datac(!Xd_0__inst_mult_5_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_219 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_228 ),
	.cout(Xd_0__inst_mult_5_229 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_303 ),
	.datab(!Xd_0__inst_mult_5_84 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_224 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_233 ),
	.cout(Xd_0__inst_mult_5_234 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_61 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[34]),
	.datac(!Xd_0__inst_mult_4_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_214 ),
	.cout(Xd_0__inst_mult_4_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_304 ),
	.datab(!Xd_0__inst_mult_4_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_219 ),
	.cout(Xd_0__inst_mult_4_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_60 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_3_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_209 ),
	.cout(Xd_0__inst_mult_3_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_299 ),
	.datab(!Xd_0__inst_mult_3_304 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_214 ),
	.cout(Xd_0__inst_mult_3_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_59 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[18]),
	.datac(!Xd_0__inst_mult_2_299 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_204 ),
	.cout(Xd_0__inst_mult_2_205 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_60 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_304 ),
	.datab(!Xd_0__inst_mult_2_309 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_209 ),
	.cout(Xd_0__inst_mult_2_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_60 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[10]),
	.datac(!Xd_0__inst_mult_1_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_209 ),
	.cout(Xd_0__inst_mult_1_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_299 ),
	.datab(!Xd_0__inst_mult_1_304 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_214 ),
	.cout(Xd_0__inst_mult_1_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_60 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_304 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_209 ),
	.cout(Xd_0__inst_mult_0_210 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_309 ),
	.datab(!Xd_0__inst_mult_0_314 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_214 ),
	.cout(Xd_0__inst_mult_0_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_214 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_314 ),
	.datab(!Xd_0__inst_mult_31_319 ),
	.datac(!din_a[253]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_219 ),
	.cout(Xd_0__inst_mult_31_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_64 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_229 ),
	.cout(Xd_0__inst_mult_30_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_269 ),
	.datab(!Xd_0__inst_mult_30_324 ),
	.datac(!din_a[245]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_234 ),
	.cout(Xd_0__inst_mult_30_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_214 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_309 ),
	.datab(!Xd_0__inst_mult_29_314 ),
	.datac(!din_a[237]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_219 ),
	.cout(Xd_0__inst_mult_29_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_62 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_219 ),
	.cout(Xd_0__inst_mult_28_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_314 ),
	.datab(!Xd_0__inst_mult_28_319 ),
	.datac(!din_a[229]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_224 ),
	.cout(Xd_0__inst_mult_28_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_214 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_309 ),
	.datab(!Xd_0__inst_mult_27_314 ),
	.datac(!din_a[221]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_219 ),
	.cout(Xd_0__inst_mult_27_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_64 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_229 ),
	.cout(Xd_0__inst_mult_26_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_269 ),
	.datab(!Xd_0__inst_mult_26_324 ),
	.datac(!din_a[213]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_234 ),
	.cout(Xd_0__inst_mult_26_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_63 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_224 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_249 ),
	.datab(!Xd_0__inst_mult_25_324 ),
	.datac(!din_a[205]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_229 ),
	.cout(Xd_0__inst_mult_25_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_63 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_224 ),
	.cout(Xd_0__inst_mult_24_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_259 ),
	.datab(!Xd_0__inst_mult_24_324 ),
	.datac(!din_a[197]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_229 ),
	.cout(Xd_0__inst_mult_24_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_234 ),
	.cout(Xd_0__inst_mult_23_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_66 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_259 ),
	.datab(!Xd_0__inst_mult_23_324 ),
	.datac(!din_a[189]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_239 ),
	.cout(Xd_0__inst_mult_23_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_234 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_66 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_259 ),
	.datab(!Xd_0__inst_mult_22_324 ),
	.datac(!din_a[181]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_239 ),
	.cout(Xd_0__inst_mult_22_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_234 ),
	.cout(Xd_0__inst_mult_21_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_66 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_259 ),
	.datab(!Xd_0__inst_mult_21_324 ),
	.datac(!din_a[173]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_239 ),
	.cout(Xd_0__inst_mult_21_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_239 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_248 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_69 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_273 ),
	.datab(!Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[165]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_253 ),
	.cout(Xd_0__inst_mult_20_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_239 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_248 ),
	.cout(Xd_0__inst_mult_19_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_69 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_273 ),
	.datab(!Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[157]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_253 ),
	.cout(Xd_0__inst_mult_19_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_239 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_248 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_69 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_273 ),
	.datab(!Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[149]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_253 ),
	.cout(Xd_0__inst_mult_18_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_239 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_248 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_69 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_273 ),
	.datab(!Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[141]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_253 ),
	.cout(Xd_0__inst_mult_17_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_239 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_248 ),
	.cout(Xd_0__inst_mult_16_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_69 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_273 ),
	.datab(!Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[133]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_253 ),
	.cout(Xd_0__inst_mult_16_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_67 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_243 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_318 ),
	.datab(!Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[125]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_239 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_248 ),
	.cout(Xd_0__inst_mult_15_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_238 ),
	.cout(Xd_0__inst_mult_14_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_308 ),
	.datab(!Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[117]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_243 ),
	.cout(Xd_0__inst_mult_14_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_238 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_313 ),
	.datab(!Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[109]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_243 ),
	.cout(Xd_0__inst_mult_13_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_238 ),
	.cout(Xd_0__inst_mult_12_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_308 ),
	.datab(!Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[101]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_243 ),
	.cout(Xd_0__inst_mult_12_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_238 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_313 ),
	.datab(!Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[93]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_243 ),
	.cout(Xd_0__inst_mult_11_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_238 ),
	.cout(Xd_0__inst_mult_10_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_313 ),
	.datab(!Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[85]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_243 ),
	.cout(Xd_0__inst_mult_10_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_238 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_308 ),
	.datab(!Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[77]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_243 ),
	.cout(Xd_0__inst_mult_9_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_238 ),
	.cout(Xd_0__inst_mult_8_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_313 ),
	.datab(!Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[69]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_243 ),
	.cout(Xd_0__inst_mult_8_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_238 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_308 ),
	.datab(!Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[61]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_243 ),
	.cout(Xd_0__inst_mult_7_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_238 ),
	.cout(Xd_0__inst_mult_6_239 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_313 ),
	.datab(!Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[53]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_243 ),
	.cout(Xd_0__inst_mult_6_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_229 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_238 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_308 ),
	.datab(!Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ),
	.datac(!din_a[45]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_234 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_243 ),
	.cout(Xd_0__inst_mult_5_244 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_63 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_224 ),
	.cout(Xd_0__inst_mult_4_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_314 ),
	.datab(!Xd_0__inst_mult_4_319 ),
	.datac(!din_a[37]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_229 ),
	.cout(Xd_0__inst_mult_4_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_62 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_219 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_309 ),
	.datab(!Xd_0__inst_mult_3_314 ),
	.datac(!din_a[29]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_224 ),
	.cout(Xd_0__inst_mult_3_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_205 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_214 ),
	.cout(Xd_0__inst_mult_2_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_62 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_314 ),
	.datab(!Xd_0__inst_mult_2_319 ),
	.datac(!din_a[21]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_219 ),
	.cout(Xd_0__inst_mult_2_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_62 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_219 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_309 ),
	.datab(!Xd_0__inst_mult_1_314 ),
	.datac(!din_a[13]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_224 ),
	.cout(Xd_0__inst_mult_1_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_62 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_210 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_219 ),
	.cout(Xd_0__inst_mult_0_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_319 ),
	.datab(!Xd_0__inst_mult_0_324 ),
	.datac(!din_a[5]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_224 ),
	.cout(Xd_0__inst_mult_0_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_314 ),
	.datab(!Xd_0__inst_mult_31_319 ),
	.datac(!Xd_0__inst_mult_31_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_224 ),
	.cout(Xd_0__inst_mult_31_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_28 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[252]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_28_sumout ),
	.cout(Xd_0__inst_mult_31_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_66 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_269 ),
	.datab(!Xd_0__inst_mult_30_324 ),
	.datac(!Xd_0__inst_mult_30_174 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_239 ),
	.cout(Xd_0__inst_mult_30_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_28 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[244]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_28_sumout ),
	.cout(Xd_0__inst_mult_30_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_309 ),
	.datab(!Xd_0__inst_mult_29_314 ),
	.datac(!Xd_0__inst_mult_29_319 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_224 ),
	.cout(Xd_0__inst_mult_29_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_28 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[236]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_28_sumout ),
	.cout(Xd_0__inst_mult_29_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_314 ),
	.datab(!Xd_0__inst_mult_28_319 ),
	.datac(!Xd_0__inst_mult_28_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_229 ),
	.cout(Xd_0__inst_mult_28_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_28 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[228]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_28_sumout ),
	.cout(Xd_0__inst_mult_28_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_309 ),
	.datab(!Xd_0__inst_mult_27_314 ),
	.datac(!Xd_0__inst_mult_27_319 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_224 ),
	.cout(Xd_0__inst_mult_27_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_28 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[220]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_28_sumout ),
	.cout(Xd_0__inst_mult_27_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_66 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_269 ),
	.datab(!Xd_0__inst_mult_26_324 ),
	.datac(!Xd_0__inst_mult_26_174 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_239 ),
	.cout(Xd_0__inst_mult_26_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_28 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[212]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_28_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_249 ),
	.datab(!Xd_0__inst_mult_25_324 ),
	.datac(!Xd_0__inst_mult_25_159 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_234 ),
	.cout(Xd_0__inst_mult_25_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_28 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[204]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_28_sumout ),
	.cout(Xd_0__inst_mult_25_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_259 ),
	.datab(!Xd_0__inst_mult_24_324 ),
	.datac(!Xd_0__inst_mult_24_169 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_234 ),
	.cout(Xd_0__inst_mult_24_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_28 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[196]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_28_sumout ),
	.cout(Xd_0__inst_mult_24_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_259 ),
	.datab(!Xd_0__inst_mult_23_324 ),
	.datac(!Xd_0__inst_mult_23_164 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_244 ),
	.cout(Xd_0__inst_mult_23_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_33 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[188]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_33_sumout ),
	.cout(Xd_0__inst_mult_23_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_259 ),
	.datab(!Xd_0__inst_mult_22_324 ),
	.datac(!Xd_0__inst_mult_22_164 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_244 ),
	.cout(Xd_0__inst_mult_22_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_33 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_33_sumout ),
	.cout(Xd_0__inst_mult_22_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_67 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_259 ),
	.datab(!Xd_0__inst_mult_21_324 ),
	.datac(!Xd_0__inst_mult_21_164 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_244 ),
	.cout(Xd_0__inst_mult_21_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_28 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[172]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_28_sumout ),
	.cout(Xd_0__inst_mult_21_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_70 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_273 ),
	.datab(!Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_20_178 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_258 ),
	.cout(Xd_0__inst_mult_20_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_23 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[164]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_23_sumout ),
	.cout(Xd_0__inst_mult_20_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_70 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_273 ),
	.datab(!Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_19_178 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_258 ),
	.cout(Xd_0__inst_mult_19_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_23 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_23_sumout ),
	.cout(Xd_0__inst_mult_19_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_70 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_273 ),
	.datab(!Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_18_178 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_258 ),
	.cout(Xd_0__inst_mult_18_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_23 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[148]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_23_sumout ),
	.cout(Xd_0__inst_mult_18_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_70 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_273 ),
	.datab(!Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_17_178 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_258 ),
	.cout(Xd_0__inst_mult_17_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_23 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[140]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_23_sumout ),
	.cout(Xd_0__inst_mult_17_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_70 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_273 ),
	.datab(!Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_16_178 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_258 ),
	.cout(Xd_0__inst_mult_16_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_69 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_318 ),
	.datab(!Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_15_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_253 ),
	.cout(Xd_0__inst_mult_15_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_23 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[124]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_23_sumout ),
	.cout(Xd_0__inst_mult_15_24 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_308 ),
	.datab(!Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_14_313 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_248 ),
	.cout(Xd_0__inst_mult_14_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_28 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[116]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_28_sumout ),
	.cout(Xd_0__inst_mult_14_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_313 ),
	.datab(!Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_13_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_248 ),
	.cout(Xd_0__inst_mult_13_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_28 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[108]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_28_sumout ),
	.cout(Xd_0__inst_mult_13_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_308 ),
	.datab(!Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_12_313 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_248 ),
	.cout(Xd_0__inst_mult_12_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_28 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[100]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_28_sumout ),
	.cout(Xd_0__inst_mult_12_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_313 ),
	.datab(!Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_11_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_248 ),
	.cout(Xd_0__inst_mult_11_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_28 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_28_sumout ),
	.cout(Xd_0__inst_mult_11_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_313 ),
	.datab(!Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_10_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_248 ),
	.cout(Xd_0__inst_mult_10_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_33 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_33_sumout ),
	.cout(Xd_0__inst_mult_10_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_308 ),
	.datab(!Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_9_313 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_248 ),
	.cout(Xd_0__inst_mult_9_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_28 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[76]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_28_sumout ),
	.cout(Xd_0__inst_mult_9_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_313 ),
	.datab(!Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_8_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_248 ),
	.cout(Xd_0__inst_mult_8_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_28 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_28_sumout ),
	.cout(Xd_0__inst_mult_8_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_308 ),
	.datab(!Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_7_313 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_248 ),
	.cout(Xd_0__inst_mult_7_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_28 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_28_sumout ),
	.cout(Xd_0__inst_mult_7_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_313 ),
	.datab(!Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_6_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_248 ),
	.cout(Xd_0__inst_mult_6_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_28 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[52]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_28_sumout ),
	.cout(Xd_0__inst_mult_6_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_68 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_308 ),
	.datab(!Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ),
	.datac(!Xd_0__inst_mult_5_313 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_244 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_248 ),
	.cout(Xd_0__inst_mult_5_249 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_33 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_33_sumout ),
	.cout(Xd_0__inst_mult_5_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_65 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_314 ),
	.datab(!Xd_0__inst_mult_4_319 ),
	.datac(!Xd_0__inst_mult_4_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_234 ),
	.cout(Xd_0__inst_mult_4_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_28 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_28_sumout ),
	.cout(Xd_0__inst_mult_4_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_309 ),
	.datab(!Xd_0__inst_mult_3_314 ),
	.datac(!Xd_0__inst_mult_3_319 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_229 ),
	.cout(Xd_0__inst_mult_3_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_28 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_28_sumout ),
	.cout(Xd_0__inst_mult_3_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_63 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_314 ),
	.datab(!Xd_0__inst_mult_2_319 ),
	.datac(!Xd_0__inst_mult_2_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_224 ),
	.cout(Xd_0__inst_mult_2_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_28 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_28_sumout ),
	.cout(Xd_0__inst_mult_2_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_309 ),
	.datab(!Xd_0__inst_mult_1_314 ),
	.datac(!Xd_0__inst_mult_1_319 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_229 ),
	.cout(Xd_0__inst_mult_1_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_28 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_28_sumout ),
	.cout(Xd_0__inst_mult_1_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_64 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_319 ),
	.datab(!Xd_0__inst_mult_0_324 ),
	.datac(!Xd_0__inst_mult_0_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_229 ),
	.cout(Xd_0__inst_mult_0_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_28 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_24 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_28_sumout ),
	.cout(Xd_0__inst_mult_0_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_64 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_31_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_229 ),
	.cout(Xd_0__inst_mult_31_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_67 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[246]),
	.datac(!Xd_0__inst_mult_30_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_244 ),
	.cout(Xd_0__inst_mult_30_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_64 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[238]),
	.datac(!Xd_0__inst_mult_29_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_229 ),
	.cout(Xd_0__inst_mult_29_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_65 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_28_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_234 ),
	.cout(Xd_0__inst_mult_28_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_64 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[222]),
	.datac(!Xd_0__inst_mult_27_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_229 ),
	.cout(Xd_0__inst_mult_27_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_67 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[214]),
	.datac(!Xd_0__inst_mult_26_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_244 ),
	.cout(Xd_0__inst_mult_26_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_66 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_25_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_239 ),
	.cout(Xd_0__inst_mult_25_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_66 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[198]),
	.datac(!Xd_0__inst_mult_24_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_239 ),
	.cout(Xd_0__inst_mult_24_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_68 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[190]),
	.datac(!Xd_0__inst_mult_23_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_249 ),
	.cout(Xd_0__inst_mult_23_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_68 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_22_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_249 ),
	.cout(Xd_0__inst_mult_22_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_68 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[174]),
	.datac(!Xd_0__inst_mult_21_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_249 ),
	.cout(Xd_0__inst_mult_21_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_71 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[166]),
	.datac(!Xd_0__inst_mult_20_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_259 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_263 ),
	.cout(Xd_0__inst_mult_20_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_28 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[165]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_28_sumout ),
	.cout(Xd_0__inst_mult_20_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_71 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_19_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_259 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_263 ),
	.cout(Xd_0__inst_mult_19_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_28 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[157]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_28_sumout ),
	.cout(Xd_0__inst_mult_19_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_71 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[150]),
	.datac(!Xd_0__inst_mult_18_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_259 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_263 ),
	.cout(Xd_0__inst_mult_18_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_28 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[149]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_29 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_28_sumout ),
	.cout(Xd_0__inst_mult_18_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_71 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[142]),
	.datac(!Xd_0__inst_mult_17_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_259 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_263 ),
	.cout(Xd_0__inst_mult_17_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_28 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[141]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_28_sumout ),
	.cout(Xd_0__inst_mult_17_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_71 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_16_163 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_259 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_263 ),
	.cout(Xd_0__inst_mult_16_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_70 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[126]),
	.datac(!Xd_0__inst_mult_15_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_258 ),
	.cout(Xd_0__inst_mult_15_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_28 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[125]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_28_sumout ),
	.cout(Xd_0__inst_mult_15_29 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_69 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[118]),
	.datac(!Xd_0__inst_mult_14_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_253 ),
	.cout(Xd_0__inst_mult_14_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_69 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_13_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_253 ),
	.cout(Xd_0__inst_mult_13_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_69 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[102]),
	.datac(!Xd_0__inst_mult_12_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_253 ),
	.cout(Xd_0__inst_mult_12_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_69 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[94]),
	.datac(!Xd_0__inst_mult_11_278 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_253 ),
	.cout(Xd_0__inst_mult_11_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_69 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_10_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_253 ),
	.cout(Xd_0__inst_mult_10_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_69 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[78]),
	.datac(!Xd_0__inst_mult_9_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_253 ),
	.cout(Xd_0__inst_mult_9_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_69 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[70]),
	.datac(!Xd_0__inst_mult_8_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_253 ),
	.cout(Xd_0__inst_mult_8_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_69 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_7_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_253 ),
	.cout(Xd_0__inst_mult_7_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_69 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[54]),
	.datac(!Xd_0__inst_mult_6_283 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_253 ),
	.cout(Xd_0__inst_mult_6_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_69 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[46]),
	.datac(!Xd_0__inst_mult_5_318 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_249 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_253 ),
	.cout(Xd_0__inst_mult_5_254 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_66 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_4_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_239 ),
	.cout(Xd_0__inst_mult_4_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_65 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[30]),
	.datac(!Xd_0__inst_mult_3_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_234 ),
	.cout(Xd_0__inst_mult_3_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_64 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[22]),
	.datac(!Xd_0__inst_mult_2_254 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_229 ),
	.cout(Xd_0__inst_mult_2_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_65 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_234 ),
	.cout(Xd_0__inst_mult_1_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_65 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[6]),
	.datac(!Xd_0__inst_mult_0_154 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_234 ),
	.cout(Xd_0__inst_mult_0_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_234 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_33 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[254]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_33_sumout ),
	.cout(Xd_0__inst_mult_31_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_249 ),
	.cout(Xd_0__inst_mult_30_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_33 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[246]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_33_sumout ),
	.cout(Xd_0__inst_mult_30_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_234 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_33 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[238]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_33_sumout ),
	.cout(Xd_0__inst_mult_29_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_239 ),
	.cout(Xd_0__inst_mult_28_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_33 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[230]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_33_sumout ),
	.cout(Xd_0__inst_mult_28_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_234 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_33 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[222]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_33_sumout ),
	.cout(Xd_0__inst_mult_27_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_68 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_249 ),
	.cout(Xd_0__inst_mult_26_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_33 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[214]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_33_sumout ),
	.cout(Xd_0__inst_mult_26_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_67 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_244 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_33 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[206]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_33_sumout ),
	.cout(Xd_0__inst_mult_25_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_67 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_244 ),
	.cout(Xd_0__inst_mult_24_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_33 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[198]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_33_sumout ),
	.cout(Xd_0__inst_mult_24_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_69 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_254 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_69 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_254 ),
	.cout(Xd_0__inst_mult_22_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_69 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_254 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_33 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[174]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_33_sumout ),
	.cout(Xd_0__inst_mult_21_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_72 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_268 ),
	.cout(Xd_0__inst_mult_20_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_33 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_33_sumout ),
	.cout(Xd_0__inst_mult_20_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_72 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_268 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_33 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[158]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_33_sumout ),
	.cout(Xd_0__inst_mult_19_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_72 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_268 ),
	.cout(Xd_0__inst_mult_18_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_33 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[150]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_33_sumout ),
	.cout(Xd_0__inst_mult_18_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_72 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_268 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_33 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_33_sumout ),
	.cout(Xd_0__inst_mult_17_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_72 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_268 ),
	.cout(Xd_0__inst_mult_16_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_33 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[134]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_33_sumout ),
	.cout(Xd_0__inst_mult_16_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_259 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_263 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_33 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[126]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_33_sumout ),
	.cout(Xd_0__inst_mult_15_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_258 ),
	.cout(Xd_0__inst_mult_14_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_33 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_33_sumout ),
	.cout(Xd_0__inst_mult_14_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_258 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_33 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[110]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_33_sumout ),
	.cout(Xd_0__inst_mult_13_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_258 ),
	.cout(Xd_0__inst_mult_12_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_33 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[102]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_33_sumout ),
	.cout(Xd_0__inst_mult_12_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_258 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_33 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_33_sumout ),
	.cout(Xd_0__inst_mult_11_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_258 ),
	.cout(Xd_0__inst_mult_10_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_258 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_33 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[78]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_33_sumout ),
	.cout(Xd_0__inst_mult_9_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_258 ),
	.cout(Xd_0__inst_mult_8_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_33 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_33_sumout ),
	.cout(Xd_0__inst_mult_8_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_258 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_33 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[62]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_33_sumout ),
	.cout(Xd_0__inst_mult_7_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_258 ),
	.cout(Xd_0__inst_mult_6_259 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_33 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_33_sumout ),
	.cout(Xd_0__inst_mult_6_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_70 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_254 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_258 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_67 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_244 ),
	.cout(Xd_0__inst_mult_4_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_33 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[38]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_33_sumout ),
	.cout(Xd_0__inst_mult_4_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_239 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_33 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_33_sumout ),
	.cout(Xd_0__inst_mult_3_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_65 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_234 ),
	.cout(Xd_0__inst_mult_2_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_33 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_33_sumout ),
	.cout(Xd_0__inst_mult_2_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_239 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_33 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[14]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_33_sumout ),
	.cout(Xd_0__inst_mult_1_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_239 ),
	.cout(Xd_0__inst_mult_0_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_33 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_34 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_33_sumout ),
	.cout(Xd_0__inst_mult_0_34 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_72 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[125]),
	.datac(!din_a[124]),
	.datad(!din_b[126]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_268 ),
	.cout(Xd_0__inst_mult_15_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_69 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[242]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_254 ),
	.cout(Xd_0__inst_mult_30_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_67 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[226]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_244 ),
	.cout(Xd_0__inst_mult_28_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_67 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[5]),
	.datac(!din_a[4]),
	.datad(!din_b[6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_244 ),
	.cout(Xd_0__inst_mult_0_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_69 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[210]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_254 ),
	.cout(Xd_0__inst_mult_26_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_67 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[26]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_244 ),
	.cout(Xd_0__inst_mult_3_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_67 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_244 ),
	.cout(Xd_0__inst_mult_1_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_66 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[249]),
	.datac(!din_a[249]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_239 ),
	.cout(Xd_0__inst_mult_31_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_31_67 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[249]),
	.datac(!din_a[249]),
	.datad(!din_b[248]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_230 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_70 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[189]),
	.datac(!din_a[187]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_259 ),
	.cout(Xd_0__inst_mult_23_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_70 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[241]),
	.datac(!din_a[241]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_259 ),
	.cout(Xd_0__inst_mult_30_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_30_71 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[241]),
	.datac(!din_a[241]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_152 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_70 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[181]),
	.datac(!din_a[179]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_259 ),
	.cout(Xd_0__inst_mult_22_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_66 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[233]),
	.datac(!din_a[233]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_239 ),
	.cout(Xd_0__inst_mult_29_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_29_67 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[233]),
	.datac(!din_a[233]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_220 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_70 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[173]),
	.datac(!din_a[171]),
	.datad(!din_b[174]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_259 ),
	.cout(Xd_0__inst_mult_21_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_68 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[225]),
	.datac(!din_a[225]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_249 ),
	.cout(Xd_0__inst_mult_28_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_28_69 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[225]),
	.datac(!din_a[225]),
	.datad(!din_b[224]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_29 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_73 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[165]),
	.datac(!din_a[163]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_273 ),
	.cout(Xd_0__inst_mult_20_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_66 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[217]),
	.datac(!din_a[217]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_239 ),
	.cout(Xd_0__inst_mult_27_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_27_67 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[217]),
	.datac(!din_a[217]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_230 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_68 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[205]),
	.datac(!din_a[203]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_249 ),
	.cout(Xd_0__inst_mult_25_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_70 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[209]),
	.datac(!din_a[209]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_259 ),
	.cout(Xd_0__inst_mult_26_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_26_71 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[209]),
	.datac(!din_a[209]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_29 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_73 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[157]),
	.datac(!din_a[155]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_273 ),
	.cout(Xd_0__inst_mult_19_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_69 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[201]),
	.datac(!din_a[201]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_254 ),
	.cout(Xd_0__inst_mult_25_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_25_70 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[201]),
	.datac(!din_a[201]),
	.datad(!din_b[200]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_235 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_73 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[149]),
	.datac(!din_a[147]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_273 ),
	.cout(Xd_0__inst_mult_18_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_68 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[193]),
	.datac(!din_a[193]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_249 ),
	.cout(Xd_0__inst_mult_24_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_24_69 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[193]),
	.datac(!din_a[193]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_34 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_73 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[141]),
	.datac(!din_a[139]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_273 ),
	.cout(Xd_0__inst_mult_17_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_71 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[185]),
	.datac(!din_a[185]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_264 ),
	.cout(Xd_0__inst_mult_23_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_23_72 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[185]),
	.datac(!din_a[185]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_34 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_70 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[197]),
	.datac(!din_a[195]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_259 ),
	.cout(Xd_0__inst_mult_24_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_71 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[177]),
	.datac(!din_a[177]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_264 ),
	.cout(Xd_0__inst_mult_22_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_22_72 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[177]),
	.datac(!din_a[177]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_235 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_68 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[33]),
	.datac(!din_a[36]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_249 ),
	.cout(Xd_0__inst_mult_4_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_71 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[169]),
	.datac(!din_a[169]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_264 ),
	.cout(Xd_0__inst_mult_21_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_21_72 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[169]),
	.datac(!din_a[169]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_29 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_72 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[213]),
	.datac(!din_a[211]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_269 ),
	.cout(Xd_0__inst_mult_26_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_74 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[161]),
	.datac(!din_a[161]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_278 ),
	.cout(Xd_0__inst_mult_20_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_20_75 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[161]),
	.datac(!din_a[161]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_249 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_73 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[133]),
	.datac(!din_a[131]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_273 ),
	.cout(Xd_0__inst_mult_16_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_74 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[153]),
	.datac(!din_a[153]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_278 ),
	.cout(Xd_0__inst_mult_19_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_19_75 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[153]),
	.datac(!din_a[153]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_24 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_71 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[97]),
	.datac(!din_a[100]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_263 ),
	.cout(Xd_0__inst_mult_12_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_74 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[145]),
	.datac(!din_a[145]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_278 ),
	.cout(Xd_0__inst_mult_18_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_18_75 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[145]),
	.datac(!din_a[145]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_225 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_73 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[185]),
	.datac(!din_a[188]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_274 ),
	.cout(Xd_0__inst_mult_23_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_74 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[137]),
	.datac(!din_a[137]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_278 ),
	.cout(Xd_0__inst_mult_17_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_17_75 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[137]),
	.datac(!din_a[137]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_249 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_71 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[41]),
	.datac(!din_a[44]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_263 ),
	.cout(Xd_0__inst_mult_5_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_74 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[129]),
	.datac(!din_a[129]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_278 ),
	.cout(Xd_0__inst_mult_16_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_16_75 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[129]),
	.datac(!din_a[129]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_132 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_71 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[49]),
	.datac(!din_a[52]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_263 ),
	.cout(Xd_0__inst_mult_6_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_73 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[121]),
	.datac(!din_a[121]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_273 ),
	.cout(Xd_0__inst_mult_15_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_15_74 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[121]),
	.datac(!din_a[121]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_239 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_71 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[57]),
	.datac(!din_a[60]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_263 ),
	.cout(Xd_0__inst_mult_7_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_71 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[113]),
	.datac(!din_a[113]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_263 ),
	.cout(Xd_0__inst_mult_14_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_14_72 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[113]),
	.datac(!din_a[113]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_320 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_71 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[65]),
	.datac(!din_a[68]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_263 ),
	.cout(Xd_0__inst_mult_8_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_71 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[105]),
	.datac(!din_a[105]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_263 ),
	.cout(Xd_0__inst_mult_13_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_13_72 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[105]),
	.datac(!din_a[105]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_239 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_71 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[73]),
	.datac(!din_a[76]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_263 ),
	.cout(Xd_0__inst_mult_9_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_72 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[97]),
	.datac(!din_a[97]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_268 ),
	.cout(Xd_0__inst_mult_12_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_12_73 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[97]),
	.datac(!din_a[97]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_315 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_76 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[153]),
	.datac(!din_a[156]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_288 ),
	.cout(Xd_0__inst_mult_19_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_71 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[89]),
	.datac(!din_a[89]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_263 ),
	.cout(Xd_0__inst_mult_11_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_11_72 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[89]),
	.datac(!din_a[89]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_239 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_71 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[81]),
	.datac(!din_a[84]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_263 ),
	.cout(Xd_0__inst_mult_10_264 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_72 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[81]),
	.datac(!din_a[81]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_268 ),
	.cout(Xd_0__inst_mult_10_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_10_73 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[81]),
	.datac(!din_a[81]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_320 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_73 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[89]),
	.datac(!din_a[92]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_273 ),
	.cout(Xd_0__inst_mult_11_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_72 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[73]),
	.datac(!din_a[73]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_268 ),
	.cout(Xd_0__inst_mult_9_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_9_73 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[73]),
	.datac(!din_a[73]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_239 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_73 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[105]),
	.datac(!din_a[108]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_273 ),
	.cout(Xd_0__inst_mult_13_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_72 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[65]),
	.datac(!din_a[65]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_268 ),
	.cout(Xd_0__inst_mult_8_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_8_73 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[65]),
	.datac(!din_a[65]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_315 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_73 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[113]),
	.datac(!din_a[116]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_273 ),
	.cout(Xd_0__inst_mult_14_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_72 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[57]),
	.datac(!din_a[57]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_268 ),
	.cout(Xd_0__inst_mult_7_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_7_73 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[57]),
	.datac(!din_a[57]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_239 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_75 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[121]),
	.datac(!din_a[124]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_283 ),
	.cout(Xd_0__inst_mult_15_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_72 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[49]),
	.datac(!din_a[49]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_268 ),
	.cout(Xd_0__inst_mult_6_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_6_73 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[49]),
	.datac(!din_a[49]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_76 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[129]),
	.datac(!din_a[132]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_288 ),
	.cout(Xd_0__inst_mult_16_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_72 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[41]),
	.datac(!din_a[41]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_159 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_268 ),
	.cout(Xd_0__inst_mult_5_269 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_5_73 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[41]),
	.datac(!din_a[41]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_225 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_274 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_76 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[137]),
	.datac(!din_a[140]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_288 ),
	.cout(Xd_0__inst_mult_17_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_69 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[33]),
	.datac(!din_a[33]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_254 ),
	.cout(Xd_0__inst_mult_4_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_4_70 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[33]),
	.datac(!din_a[33]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_315 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_76 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[145]),
	.datac(!din_a[148]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_288 ),
	.cout(Xd_0__inst_mult_18_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_68 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[25]),
	.datac(!din_a[25]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_249 ),
	.cout(Xd_0__inst_mult_3_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_3_69 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[25]),
	.datac(!din_a[25]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_215 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_72 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[245]),
	.datac(!din_a[243]),
	.datad(!din_b[246]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_269 ),
	.cout(Xd_0__inst_mult_30_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_66 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[17]),
	.datac(!din_a[17]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_239 ),
	.cout(Xd_0__inst_mult_2_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_2_67 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[17]),
	.datac(!din_a[17]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_320 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_76 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[161]),
	.datac(!din_a[164]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_288 ),
	.cout(Xd_0__inst_mult_20_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_68 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[9]),
	.datac(!din_a[9]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_249 ),
	.cout(Xd_0__inst_mult_1_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_1_69 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[9]),
	.datac(!din_a[9]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_220 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_73 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[169]),
	.datac(!din_a[172]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_274 ),
	.cout(Xd_0__inst_mult_21_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_68 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[1]),
	.datac(!din_a[1]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_150 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_249 ),
	.cout(Xd_0__inst_mult_0_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_0_69 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[1]),
	.datac(!din_a[1]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_73 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[177]),
	.datac(!din_a[180]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_274 ),
	.cout(Xd_0__inst_mult_22_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_68 (
// Equation(s):

	.dataa(!din_a[251]),
	.datab(!din_b[249]),
	.datac(!din_a[250]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_249 ),
	.cout(Xd_0__inst_mult_31_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_73 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[241]),
	.datac(!din_a[242]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_274 ),
	.cout(Xd_0__inst_mult_30_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_68 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[233]),
	.datac(!din_a[234]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_249 ),
	.cout(Xd_0__inst_mult_29_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_69 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_254 ),
	.cout(Xd_0__inst_mult_31_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_70 (
// Equation(s):

	.dataa(!din_a[227]),
	.datab(!din_b[225]),
	.datac(!din_a[226]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_259 ),
	.cout(Xd_0__inst_mult_28_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_68 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[217]),
	.datac(!din_a[218]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_249 ),
	.cout(Xd_0__inst_mult_27_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_264 ),
	.cout(Xd_0__inst_mult_28_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_73 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[209]),
	.datac(!din_a[210]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_274 ),
	.cout(Xd_0__inst_mult_26_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_71 (
// Equation(s):

	.dataa(!din_a[203]),
	.datab(!din_b[201]),
	.datac(!din_a[202]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_264 ),
	.cout(Xd_0__inst_mult_25_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_71 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[193]),
	.datac(!din_a[194]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_264 ),
	.cout(Xd_0__inst_mult_24_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_74 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[185]),
	.datac(!din_a[186]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_279 ),
	.cout(Xd_0__inst_mult_23_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_74 (
// Equation(s):

	.dataa(!din_a[179]),
	.datab(!din_b[177]),
	.datac(!din_a[178]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_279 ),
	.cout(Xd_0__inst_mult_22_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_74 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[169]),
	.datac(!din_a[170]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_279 ),
	.cout(Xd_0__inst_mult_21_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_77 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[161]),
	.datac(!din_a[162]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_293 ),
	.cout(Xd_0__inst_mult_20_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_77 (
// Equation(s):

	.dataa(!din_a[155]),
	.datab(!din_b[153]),
	.datac(!din_a[154]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_293 ),
	.cout(Xd_0__inst_mult_19_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_77 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[145]),
	.datac(!din_a[146]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_293 ),
	.cout(Xd_0__inst_mult_18_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_77 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[137]),
	.datac(!din_a[138]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_293 ),
	.cout(Xd_0__inst_mult_17_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_77 (
// Equation(s):

	.dataa(!din_a[131]),
	.datab(!din_b[129]),
	.datac(!din_a[130]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_293 ),
	.cout(Xd_0__inst_mult_16_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_76 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[121]),
	.datac(!din_a[122]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_274 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_288 ),
	.cout(Xd_0__inst_mult_15_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_74 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[113]),
	.datac(!din_a[114]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_278 ),
	.cout(Xd_0__inst_mult_14_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_74 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_278 ),
	.cout(Xd_0__inst_mult_13_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_75 (
// Equation(s):

	.dataa(!din_a[107]),
	.datab(!din_b[105]),
	.datac(!din_a[106]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_283 ),
	.cout(Xd_0__inst_mult_13_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_74 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[97]),
	.datac(!din_a[98]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_278 ),
	.cout(Xd_0__inst_mult_12_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_74 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_278 ),
	.cout(Xd_0__inst_mult_11_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_75 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[89]),
	.datac(!din_a[90]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_264 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_283 ),
	.cout(Xd_0__inst_mult_11_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_74 (
// Equation(s):

	.dataa(!din_a[83]),
	.datab(!din_b[81]),
	.datac(!din_a[82]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_278 ),
	.cout(Xd_0__inst_mult_10_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_74 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_278 ),
	.cout(Xd_0__inst_mult_9_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_75 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_283 ),
	.cout(Xd_0__inst_mult_10_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_74 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[65]),
	.datac(!din_a[66]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_278 ),
	.cout(Xd_0__inst_mult_8_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_74 (
// Equation(s):

	.dataa(!din_a[59]),
	.datab(!din_b[57]),
	.datac(!din_a[58]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_278 ),
	.cout(Xd_0__inst_mult_7_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_75 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_283 ),
	.cout(Xd_0__inst_mult_8_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_74 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[49]),
	.datac(!din_a[50]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_278 ),
	.cout(Xd_0__inst_mult_6_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_74 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[41]),
	.datac(!din_a[42]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_269 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_278 ),
	.cout(Xd_0__inst_mult_5_279 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_75 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_319 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_283 ),
	.cout(Xd_0__inst_mult_6_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_71 (
// Equation(s):

	.dataa(!din_a[35]),
	.datab(!din_b[33]),
	.datac(!din_a[34]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_264 ),
	.cout(Xd_0__inst_mult_4_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_70 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[25]),
	.datac(!din_a[26]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_259 ),
	.cout(Xd_0__inst_mult_3_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_72 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_269 ),
	.cout(Xd_0__inst_mult_4_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_68 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[17]),
	.datac(!din_a[18]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_249 ),
	.cout(Xd_0__inst_mult_2_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_70 (
// Equation(s):

	.dataa(!din_a[11]),
	.datab(!din_b[9]),
	.datac(!din_a[10]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_259 ),
	.cout(Xd_0__inst_mult_1_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_69 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_254 ),
	.cout(Xd_0__inst_mult_2_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_70 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_259 ),
	.cout(Xd_0__inst_mult_0_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_70 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[249]),
	.datac(!din_a[251]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_259 ),
	.cout(Xd_0__inst_mult_31_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_74 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[241]),
	.datac(!din_a[243]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_279 ),
	.cout(Xd_0__inst_mult_30_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_69 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[233]),
	.datac(!din_a[235]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_254 ),
	.cout(Xd_0__inst_mult_29_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_72 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[225]),
	.datac(!din_a[227]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_269 ),
	.cout(Xd_0__inst_mult_28_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_69 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[217]),
	.datac(!din_a[219]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_254 ),
	.cout(Xd_0__inst_mult_27_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_74 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[209]),
	.datac(!din_a[211]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_279 ),
	.cout(Xd_0__inst_mult_26_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_72 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[201]),
	.datac(!din_a[203]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_269 ),
	.cout(Xd_0__inst_mult_25_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_72 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[193]),
	.datac(!din_a[195]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_269 ),
	.cout(Xd_0__inst_mult_24_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_75 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[185]),
	.datac(!din_a[187]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_284 ),
	.cout(Xd_0__inst_mult_23_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_75 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[177]),
	.datac(!din_a[179]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_284 ),
	.cout(Xd_0__inst_mult_22_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_75 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[169]),
	.datac(!din_a[171]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_284 ),
	.cout(Xd_0__inst_mult_21_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_78 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[161]),
	.datac(!din_a[163]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_298 ),
	.cout(Xd_0__inst_mult_20_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_78 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[153]),
	.datac(!din_a[155]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_298 ),
	.cout(Xd_0__inst_mult_19_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_78 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[145]),
	.datac(!din_a[147]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_298 ),
	.cout(Xd_0__inst_mult_18_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_78 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[137]),
	.datac(!din_a[139]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_298 ),
	.cout(Xd_0__inst_mult_17_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_78 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[129]),
	.datac(!din_a[131]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_298 ),
	.cout(Xd_0__inst_mult_16_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_77 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[121]),
	.datac(!din_a[123]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_293 ),
	.cout(Xd_0__inst_mult_15_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_75 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[113]),
	.datac(!din_a[115]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_283 ),
	.cout(Xd_0__inst_mult_14_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_76 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[105]),
	.datac(!din_a[107]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_288 ),
	.cout(Xd_0__inst_mult_13_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_75 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[97]),
	.datac(!din_a[99]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_283 ),
	.cout(Xd_0__inst_mult_12_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_76 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[89]),
	.datac(!din_a[91]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_284 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_288 ),
	.cout(Xd_0__inst_mult_11_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_76 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[81]),
	.datac(!din_a[83]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_288 ),
	.cout(Xd_0__inst_mult_10_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_75 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[73]),
	.datac(!din_a[75]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_283 ),
	.cout(Xd_0__inst_mult_9_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_76 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[65]),
	.datac(!din_a[67]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_288 ),
	.cout(Xd_0__inst_mult_8_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_75 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[57]),
	.datac(!din_a[59]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_283 ),
	.cout(Xd_0__inst_mult_7_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_76 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[49]),
	.datac(!din_a[51]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_288 ),
	.cout(Xd_0__inst_mult_6_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_75 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[41]),
	.datac(!din_a[43]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_279 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_283 ),
	.cout(Xd_0__inst_mult_5_284 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_73 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[33]),
	.datac(!din_a[35]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_274 ),
	.cout(Xd_0__inst_mult_4_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_71 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[25]),
	.datac(!din_a[27]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_264 ),
	.cout(Xd_0__inst_mult_3_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_70 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[17]),
	.datac(!din_a[19]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_259 ),
	.cout(Xd_0__inst_mult_2_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_71 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[9]),
	.datac(!din_a[11]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_264 ),
	.cout(Xd_0__inst_mult_1_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_71 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[1]),
	.datac(!din_a[3]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_264 ),
	.cout(Xd_0__inst_mult_0_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_71 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[249]),
	.datac(!din_a[252]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_264 ),
	.cout(Xd_0__inst_mult_31_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_72 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[254]),
	.datac(!din_a[250]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_269 ),
	.cout(Xd_0__inst_mult_31_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_73 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[253]),
	.datac(!din_a[251]),
	.datad(!din_b[251]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_274 ),
	.cout(Xd_0__inst_mult_31_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_31_74 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[252]),
	.datac(!din_a[249]),
	.datad(!din_b[251]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_269 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_75 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[241]),
	.datac(!din_a[244]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_284 ),
	.cout(Xd_0__inst_mult_30_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_76 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[246]),
	.datac(!din_a[242]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_289 ),
	.cout(Xd_0__inst_mult_30_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_77 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[245]),
	.datac(!din_a[243]),
	.datad(!din_b[243]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_294 ),
	.cout(Xd_0__inst_mult_30_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_30_78 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[244]),
	.datac(!din_a[241]),
	.datad(!din_b[243]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_112 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_70 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[233]),
	.datac(!din_a[236]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_259 ),
	.cout(Xd_0__inst_mult_29_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_71 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[238]),
	.datac(!din_a[234]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_264 ),
	.cout(Xd_0__inst_mult_29_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_72 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[237]),
	.datac(!din_a[235]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_269 ),
	.cout(Xd_0__inst_mult_29_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_29_73 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[236]),
	.datac(!din_a[233]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_250 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_73 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[225]),
	.datac(!din_a[228]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_274 ),
	.cout(Xd_0__inst_mult_28_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_74 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[230]),
	.datac(!din_a[226]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_279 ),
	.cout(Xd_0__inst_mult_28_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_75 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[229]),
	.datac(!din_a[227]),
	.datad(!din_b[227]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_284 ),
	.cout(Xd_0__inst_mult_28_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_28_76 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[228]),
	.datac(!din_a[225]),
	.datad(!din_b[227]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_92 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_70 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[217]),
	.datac(!din_a[220]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_259 ),
	.cout(Xd_0__inst_mult_27_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_71 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[222]),
	.datac(!din_a[218]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_264 ),
	.cout(Xd_0__inst_mult_27_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_72 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[221]),
	.datac(!din_a[219]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_269 ),
	.cout(Xd_0__inst_mult_27_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_27_73 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[220]),
	.datac(!din_a[217]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_240 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_75 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[209]),
	.datac(!din_a[212]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_284 ),
	.cout(Xd_0__inst_mult_26_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_76 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[214]),
	.datac(!din_a[210]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_195 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_289 ),
	.cout(Xd_0__inst_mult_26_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_77 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[213]),
	.datac(!din_a[211]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_294 ),
	.cout(Xd_0__inst_mult_26_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_26_78 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[212]),
	.datac(!din_a[209]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_77 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_73 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[201]),
	.datac(!din_a[204]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_274 ),
	.cout(Xd_0__inst_mult_25_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_74 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[206]),
	.datac(!din_a[202]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_279 ),
	.cout(Xd_0__inst_mult_25_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_75 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[205]),
	.datac(!din_a[203]),
	.datad(!din_b[203]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_284 ),
	.cout(Xd_0__inst_mult_25_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_25_76 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[204]),
	.datac(!din_a[201]),
	.datad(!din_b[203]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_250 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_73 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[193]),
	.datac(!din_a[196]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_274 ),
	.cout(Xd_0__inst_mult_24_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_74 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[198]),
	.datac(!din_a[194]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_279 ),
	.cout(Xd_0__inst_mult_24_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_75 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[197]),
	.datac(!din_a[195]),
	.datad(!din_b[195]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_284 ),
	.cout(Xd_0__inst_mult_24_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_24_76 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[196]),
	.datac(!din_a[193]),
	.datad(!din_b[195]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_52 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_76 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[190]),
	.datac(!din_a[186]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_289 ),
	.cout(Xd_0__inst_mult_23_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_77 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[189]),
	.datac(!din_a[187]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_294 ),
	.cout(Xd_0__inst_mult_23_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_23_78 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[188]),
	.datac(!din_a[185]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_245 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_76 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[182]),
	.datac(!din_a[178]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_289 ),
	.cout(Xd_0__inst_mult_22_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_77 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[181]),
	.datac(!din_a[179]),
	.datad(!din_b[179]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_294 ),
	.cout(Xd_0__inst_mult_22_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_22_78 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[180]),
	.datac(!din_a[177]),
	.datad(!din_b[179]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_32 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_76 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[174]),
	.datac(!din_a[170]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_200 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_289 ),
	.cout(Xd_0__inst_mult_21_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_77 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[173]),
	.datac(!din_a[171]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_294 ),
	.cout(Xd_0__inst_mult_21_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_21_78 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[172]),
	.datac(!din_a[169]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_255 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_79 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[166]),
	.datac(!din_a[162]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_303 ),
	.cout(Xd_0__inst_mult_20_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_20_80 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[164]),
	.datac(!din_a[161]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i21_12 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_79 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[158]),
	.datac(!din_a[154]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_303 ),
	.cout(Xd_0__inst_mult_19_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_19_80 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[156]),
	.datac(!din_a[153]),
	.datad(!din_b[155]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_269 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_79 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[150]),
	.datac(!din_a[146]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_303 ),
	.cout(Xd_0__inst_mult_18_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_18_80 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[148]),
	.datac(!din_a[145]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_34 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_79 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[142]),
	.datac(!din_a[138]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_303 ),
	.cout(Xd_0__inst_mult_17_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_17_80 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[140]),
	.datac(!din_a[137]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_269 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_79 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[134]),
	.datac(!din_a[130]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_214 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_303 ),
	.cout(Xd_0__inst_mult_16_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_16_80 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[132]),
	.datac(!din_a[129]),
	.datad(!din_b[131]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_34 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_78 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[126]),
	.datac(!din_a[122]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_209 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_298 ),
	.cout(Xd_0__inst_mult_15_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_15_79 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[124]),
	.datac(!din_a[121]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_240 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_76 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[118]),
	.datac(!din_a[114]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_288 ),
	.cout(Xd_0__inst_mult_14_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_14_77 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[116]),
	.datac(!din_a[113]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_77 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[110]),
	.datac(!din_a[106]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_293 ),
	.cout(Xd_0__inst_mult_13_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_13_78 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[108]),
	.datac(!din_a[105]),
	.datad(!din_b[107]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_259 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_76 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[102]),
	.datac(!din_a[98]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_288 ),
	.cout(Xd_0__inst_mult_12_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_12_77 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[100]),
	.datac(!din_a[97]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_320 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_77 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[94]),
	.datac(!din_a[90]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_293 ),
	.cout(Xd_0__inst_mult_11_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_11_78 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[92]),
	.datac(!din_a[89]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_259 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_77 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[86]),
	.datac(!din_a[82]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_293 ),
	.cout(Xd_0__inst_mult_10_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_10_78 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[84]),
	.datac(!din_a[81]),
	.datad(!din_b[83]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_76 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[78]),
	.datac(!din_a[74]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_288 ),
	.cout(Xd_0__inst_mult_9_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_9_77 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[76]),
	.datac(!din_a[73]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_259 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_77 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[70]),
	.datac(!din_a[66]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_293 ),
	.cout(Xd_0__inst_mult_8_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_8_78 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[68]),
	.datac(!din_a[65]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_76 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[62]),
	.datac(!din_a[58]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_288 ),
	.cout(Xd_0__inst_mult_7_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_7_77 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[60]),
	.datac(!din_a[57]),
	.datad(!din_b[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_259 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_77 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[54]),
	.datac(!din_a[50]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_293 ),
	.cout(Xd_0__inst_mult_6_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_6_78 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[52]),
	.datac(!din_a[49]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_76 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[46]),
	.datac(!din_a[42]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_204 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_288 ),
	.cout(Xd_0__inst_mult_5_289 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_5_77 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[44]),
	.datac(!din_a[41]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_259 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_294 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_74 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[38]),
	.datac(!din_a[34]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_190 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_279 ),
	.cout(Xd_0__inst_mult_4_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_75 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[37]),
	.datac(!din_a[35]),
	.datad(!din_b[35]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_284 ),
	.cout(Xd_0__inst_mult_4_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_4_76 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[36]),
	.datac(!din_a[33]),
	.datad(!din_b[35]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_72 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[25]),
	.datac(!din_a[28]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_269 ),
	.cout(Xd_0__inst_mult_3_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_73 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[30]),
	.datac(!din_a[26]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_274 ),
	.cout(Xd_0__inst_mult_3_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_74 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[29]),
	.datac(!din_a[27]),
	.datad(!din_b[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_279 ),
	.cout(Xd_0__inst_mult_3_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_3_75 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[28]),
	.datac(!din_a[25]),
	.datad(!din_b[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_245 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_71 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[17]),
	.datac(!din_a[20]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_264 ),
	.cout(Xd_0__inst_mult_2_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_72 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[22]),
	.datac(!din_a[18]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_180 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_269 ),
	.cout(Xd_0__inst_mult_2_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_73 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[21]),
	.datac(!din_a[19]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_274 ),
	.cout(Xd_0__inst_mult_2_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_2_74 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[20]),
	.datac(!din_a[17]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_315 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_72 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[9]),
	.datac(!din_a[12]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_269 ),
	.cout(Xd_0__inst_mult_1_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_73 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[14]),
	.datac(!din_a[10]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_274 ),
	.cout(Xd_0__inst_mult_1_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_74 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[13]),
	.datac(!din_a[11]),
	.datad(!din_b[11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_279 ),
	.cout(Xd_0__inst_mult_1_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_1_75 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[12]),
	.datac(!din_a[9]),
	.datad(!din_b[11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_235 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_72 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[1]),
	.datac(!din_a[4]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_269 ),
	.cout(Xd_0__inst_mult_0_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_73 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[6]),
	.datac(!din_a[2]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_185 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_274 ),
	.cout(Xd_0__inst_mult_0_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_74 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[5]),
	.datac(!din_a[3]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_279 ),
	.cout(Xd_0__inst_mult_0_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_0_75 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[4]),
	.datac(!din_a[1]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_325 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_75 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[250]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_284 ),
	.cout(Xd_0__inst_mult_31_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_76 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[254]),
	.datac(!din_a[251]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_289 ),
	.cout(Xd_0__inst_mult_31_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_77 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[253]),
	.datac(!din_a[252]),
	.datad(!din_b[251]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_294 ),
	.cout(Xd_0__inst_mult_31_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_79 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[246]),
	.datac(!din_a[243]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_304 ),
	.cout(Xd_0__inst_mult_30_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_80 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[245]),
	.datac(!din_a[244]),
	.datad(!din_b[243]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_309 ),
	.cout(Xd_0__inst_mult_30_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_74 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[234]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_279 ),
	.cout(Xd_0__inst_mult_29_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_75 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[238]),
	.datac(!din_a[235]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_284 ),
	.cout(Xd_0__inst_mult_29_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_76 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[237]),
	.datac(!din_a[236]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_289 ),
	.cout(Xd_0__inst_mult_29_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_77 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[230]),
	.datac(!din_a[227]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_294 ),
	.cout(Xd_0__inst_mult_28_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_78 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[229]),
	.datac(!din_a[228]),
	.datad(!din_b[227]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_299 ),
	.cout(Xd_0__inst_mult_28_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_74 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[218]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_279 ),
	.cout(Xd_0__inst_mult_27_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_75 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[222]),
	.datac(!din_a[219]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_284 ),
	.cout(Xd_0__inst_mult_27_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_76 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[221]),
	.datac(!din_a[220]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_289 ),
	.cout(Xd_0__inst_mult_27_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_79 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[214]),
	.datac(!din_a[211]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_304 ),
	.cout(Xd_0__inst_mult_26_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_80 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[213]),
	.datac(!din_a[212]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_309 ),
	.cout(Xd_0__inst_mult_26_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_77 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[202]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_294 ),
	.cout(Xd_0__inst_mult_25_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_78 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[206]),
	.datac(!din_a[203]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_299 ),
	.cout(Xd_0__inst_mult_25_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_79 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[205]),
	.datac(!din_a[204]),
	.datad(!din_b[203]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_304 ),
	.cout(Xd_0__inst_mult_25_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_77 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[194]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_294 ),
	.cout(Xd_0__inst_mult_24_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_78 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[198]),
	.datac(!din_a[195]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_299 ),
	.cout(Xd_0__inst_mult_24_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_79 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[197]),
	.datac(!din_a[196]),
	.datad(!din_b[195]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_304 ),
	.cout(Xd_0__inst_mult_24_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_79 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[190]),
	.datac(!din_a[187]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_304 ),
	.cout(Xd_0__inst_mult_23_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_80 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[189]),
	.datac(!din_a[188]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_309 ),
	.cout(Xd_0__inst_mult_23_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_79 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[182]),
	.datac(!din_a[179]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_304 ),
	.cout(Xd_0__inst_mult_22_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_80 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[181]),
	.datac(!din_a[180]),
	.datad(!din_b[179]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_309 ),
	.cout(Xd_0__inst_mult_22_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_79 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[174]),
	.datac(!din_a[171]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_304 ),
	.cout(Xd_0__inst_mult_21_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_80 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[173]),
	.datac(!din_a[172]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_309 ),
	.cout(Xd_0__inst_mult_21_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_81 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[166]),
	.datac(!din_a[163]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_313 ),
	.cout(Xd_0__inst_mult_20_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_81 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[158]),
	.datac(!din_a[155]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_313 ),
	.cout(Xd_0__inst_mult_19_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_81 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[150]),
	.datac(!din_a[147]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_313 ),
	.cout(Xd_0__inst_mult_18_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_81 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[142]),
	.datac(!din_a[139]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_313 ),
	.cout(Xd_0__inst_mult_17_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_81 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[134]),
	.datac(!din_a[131]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_313 ),
	.cout(Xd_0__inst_mult_16_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_80 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[126]),
	.datac(!din_a[123]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_308 ),
	.cout(Xd_0__inst_mult_15_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_78 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[118]),
	.datac(!din_a[115]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_298 ),
	.cout(Xd_0__inst_mult_14_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_79 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[110]),
	.datac(!din_a[107]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_303 ),
	.cout(Xd_0__inst_mult_13_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_78 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[102]),
	.datac(!din_a[99]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_298 ),
	.cout(Xd_0__inst_mult_12_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_79 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[94]),
	.datac(!din_a[91]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_303 ),
	.cout(Xd_0__inst_mult_11_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_79 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[86]),
	.datac(!din_a[83]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_303 ),
	.cout(Xd_0__inst_mult_10_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_78 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[78]),
	.datac(!din_a[75]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_298 ),
	.cout(Xd_0__inst_mult_9_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_79 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[70]),
	.datac(!din_a[67]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_303 ),
	.cout(Xd_0__inst_mult_8_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_78 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[62]),
	.datac(!din_a[59]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_298 ),
	.cout(Xd_0__inst_mult_7_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_79 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[54]),
	.datac(!din_a[51]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_294 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_303 ),
	.cout(Xd_0__inst_mult_6_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_78 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[46]),
	.datac(!din_a[43]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_289 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_298 ),
	.cout(Xd_0__inst_mult_5_299 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_77 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[38]),
	.datac(!din_a[35]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_294 ),
	.cout(Xd_0__inst_mult_4_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_78 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[37]),
	.datac(!din_a[36]),
	.datad(!din_b[35]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_299 ),
	.cout(Xd_0__inst_mult_4_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_76 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[30]),
	.datac(!din_a[27]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_289 ),
	.cout(Xd_0__inst_mult_3_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_77 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[29]),
	.datac(!din_a[28]),
	.datad(!din_b[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_294 ),
	.cout(Xd_0__inst_mult_3_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_75 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_284 ),
	.cout(Xd_0__inst_mult_2_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_76 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[22]),
	.datac(!din_a[19]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_289 ),
	.cout(Xd_0__inst_mult_2_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_77 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[21]),
	.datac(!din_a[20]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_294 ),
	.cout(Xd_0__inst_mult_2_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_76 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[14]),
	.datac(!din_a[11]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_289 ),
	.cout(Xd_0__inst_mult_1_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_77 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[13]),
	.datac(!din_a[12]),
	.datad(!din_b[11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_294 ),
	.cout(Xd_0__inst_mult_1_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_76 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_289 ),
	.cout(Xd_0__inst_mult_0_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_77 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[6]),
	.datac(!din_a[3]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_294 ),
	.cout(Xd_0__inst_mult_0_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_78 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[5]),
	.datac(!din_a[4]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_299 ),
	.cout(Xd_0__inst_mult_0_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_78 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_299 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_79 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[254]),
	.datac(!din_a[251]),
	.datad(!din_b[253]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_304 ),
	.cout(Xd_0__inst_mult_31_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_80 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[251]),
	.datac(!din_a[252]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_309 ),
	.cout(Xd_0__inst_mult_31_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_81 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[246]),
	.datac(!din_a[243]),
	.datad(!din_b[245]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_314 ),
	.cout(Xd_0__inst_mult_30_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_82 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[243]),
	.datac(!din_a[244]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_319 ),
	.cout(Xd_0__inst_mult_30_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_77 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_78 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[238]),
	.datac(!din_a[235]),
	.datad(!din_b[237]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_299 ),
	.cout(Xd_0__inst_mult_29_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_79 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[235]),
	.datac(!din_a[236]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_304 ),
	.cout(Xd_0__inst_mult_29_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_79 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[230]),
	.datac(!din_a[227]),
	.datad(!din_b[229]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_304 ),
	.cout(Xd_0__inst_mult_28_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_80 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[227]),
	.datac(!din_a[228]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_309 ),
	.cout(Xd_0__inst_mult_28_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_77 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_78 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[222]),
	.datac(!din_a[219]),
	.datad(!din_b[221]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_299 ),
	.cout(Xd_0__inst_mult_27_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_79 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[219]),
	.datac(!din_a[220]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_304 ),
	.cout(Xd_0__inst_mult_27_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_81 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[214]),
	.datac(!din_a[211]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_314 ),
	.cout(Xd_0__inst_mult_26_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_82 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[211]),
	.datac(!din_a[212]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_319 ),
	.cout(Xd_0__inst_mult_26_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_80 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_81 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[206]),
	.datac(!din_a[203]),
	.datad(!din_b[205]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_314 ),
	.cout(Xd_0__inst_mult_25_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_82 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[203]),
	.datac(!din_a[204]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_319 ),
	.cout(Xd_0__inst_mult_25_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_80 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_81 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[198]),
	.datac(!din_a[195]),
	.datad(!din_b[197]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_314 ),
	.cout(Xd_0__inst_mult_24_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_82 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[195]),
	.datac(!din_a[196]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_319 ),
	.cout(Xd_0__inst_mult_24_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_81 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[190]),
	.datac(!din_a[187]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_314 ),
	.cout(Xd_0__inst_mult_23_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_82 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[187]),
	.datac(!din_a[188]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_319 ),
	.cout(Xd_0__inst_mult_23_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_81 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[182]),
	.datac(!din_a[179]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_314 ),
	.cout(Xd_0__inst_mult_22_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_82 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[179]),
	.datac(!din_a[180]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_319 ),
	.cout(Xd_0__inst_mult_22_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_81 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[174]),
	.datac(!din_a[171]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_314 ),
	.cout(Xd_0__inst_mult_21_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_82 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[171]),
	.datac(!din_a[172]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_319 ),
	.cout(Xd_0__inst_mult_21_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_82 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[166]),
	.datac(!din_a[163]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_318 ),
	.cout(Xd_0__inst_mult_20_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_82 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[158]),
	.datac(!din_a[155]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_318 ),
	.cout(Xd_0__inst_mult_19_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_82 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[150]),
	.datac(!din_a[147]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_318 ),
	.cout(Xd_0__inst_mult_18_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_82 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[142]),
	.datac(!din_a[139]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_318 ),
	.cout(Xd_0__inst_mult_17_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_82 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[134]),
	.datac(!din_a[131]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_318 ),
	.cout(Xd_0__inst_mult_16_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_81 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[126]),
	.datac(!din_a[123]),
	.datad(!din_b[125]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_313 ),
	.cout(Xd_0__inst_mult_15_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_79 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[118]),
	.datac(!din_a[115]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_303 ),
	.cout(Xd_0__inst_mult_14_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_80 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[110]),
	.datac(!din_a[107]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_308 ),
	.cout(Xd_0__inst_mult_13_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_79 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[102]),
	.datac(!din_a[99]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_303 ),
	.cout(Xd_0__inst_mult_12_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_80 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[94]),
	.datac(!din_a[91]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_308 ),
	.cout(Xd_0__inst_mult_11_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_80 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[86]),
	.datac(!din_a[83]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_308 ),
	.cout(Xd_0__inst_mult_10_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_79 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[78]),
	.datac(!din_a[75]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_303 ),
	.cout(Xd_0__inst_mult_9_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_80 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[70]),
	.datac(!din_a[67]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_308 ),
	.cout(Xd_0__inst_mult_8_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_79 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[62]),
	.datac(!din_a[59]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_303 ),
	.cout(Xd_0__inst_mult_7_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_80 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[54]),
	.datac(!din_a[51]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_308 ),
	.cout(Xd_0__inst_mult_6_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_79 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[46]),
	.datac(!din_a[43]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_299 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_303 ),
	.cout(Xd_0__inst_mult_5_304 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_79 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[38]),
	.datac(!din_a[35]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_304 ),
	.cout(Xd_0__inst_mult_4_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_80 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[35]),
	.datac(!din_a[36]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_309 ),
	.cout(Xd_0__inst_mult_4_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_78 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[30]),
	.datac(!din_a[27]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_299 ),
	.cout(Xd_0__inst_mult_3_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_79 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[27]),
	.datac(!din_a[28]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_304 ),
	.cout(Xd_0__inst_mult_3_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_78 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_299 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_79 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[22]),
	.datac(!din_a[19]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_304 ),
	.cout(Xd_0__inst_mult_2_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_80 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[19]),
	.datac(!din_a[20]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_309 ),
	.cout(Xd_0__inst_mult_2_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_78 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[14]),
	.datac(!din_a[11]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_299 ),
	.cout(Xd_0__inst_mult_1_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_79 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[11]),
	.datac(!din_a[12]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_304 ),
	.cout(Xd_0__inst_mult_1_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_79 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_304 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_80 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[6]),
	.datac(!din_a[3]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_309 ),
	.cout(Xd_0__inst_mult_0_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_81 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[3]),
	.datac(!din_a[4]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_314 ),
	.cout(Xd_0__inst_mult_0_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_81 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[253]),
	.datac(!din_a[251]),
	.datad(!din_b[254]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_314 ),
	.cout(Xd_0__inst_mult_31_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_319 ),
	.cout(Xd_0__inst_mult_31_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_324 ),
	.cout(Xd_0__inst_mult_30_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_80 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[237]),
	.datac(!din_a[235]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_309 ),
	.cout(Xd_0__inst_mult_29_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_314 ),
	.cout(Xd_0__inst_mult_29_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_81 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[229]),
	.datac(!din_a[227]),
	.datad(!din_b[230]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_314 ),
	.cout(Xd_0__inst_mult_28_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_319 ),
	.cout(Xd_0__inst_mult_28_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_80 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[221]),
	.datac(!din_a[219]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_309 ),
	.cout(Xd_0__inst_mult_27_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_314 ),
	.cout(Xd_0__inst_mult_27_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_324 ),
	.cout(Xd_0__inst_mult_26_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_324 ),
	.cout(Xd_0__inst_mult_25_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_324 ),
	.cout(Xd_0__inst_mult_24_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_324 ),
	.cout(Xd_0__inst_mult_23_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_324 ),
	.cout(Xd_0__inst_mult_22_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_324 ),
	.cout(Xd_0__inst_mult_21_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_82 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[125]),
	.datac(!din_a[123]),
	.datad(!din_b[126]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_318 ),
	.cout(Xd_0__inst_mult_15_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_80 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[117]),
	.datac(!din_a[115]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_308 ),
	.cout(Xd_0__inst_mult_14_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_81 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[109]),
	.datac(!din_a[107]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_313 ),
	.cout(Xd_0__inst_mult_13_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_80 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[101]),
	.datac(!din_a[99]),
	.datad(!din_b[102]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_308 ),
	.cout(Xd_0__inst_mult_12_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_81 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[93]),
	.datac(!din_a[91]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_313 ),
	.cout(Xd_0__inst_mult_11_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_81 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[85]),
	.datac(!din_a[83]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_313 ),
	.cout(Xd_0__inst_mult_10_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_80 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[77]),
	.datac(!din_a[75]),
	.datad(!din_b[78]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_308 ),
	.cout(Xd_0__inst_mult_9_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_81 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[69]),
	.datac(!din_a[67]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_313 ),
	.cout(Xd_0__inst_mult_8_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_80 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[61]),
	.datac(!din_a[59]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_308 ),
	.cout(Xd_0__inst_mult_7_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_81 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[53]),
	.datac(!din_a[51]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_313 ),
	.cout(Xd_0__inst_mult_6_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_80 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[45]),
	.datac(!din_a[43]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_304 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_308 ),
	.cout(Xd_0__inst_mult_5_309 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_81 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[37]),
	.datac(!din_a[35]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_314 ),
	.cout(Xd_0__inst_mult_4_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_319 ),
	.cout(Xd_0__inst_mult_4_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_80 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[29]),
	.datac(!din_a[27]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_309 ),
	.cout(Xd_0__inst_mult_3_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_314 ),
	.cout(Xd_0__inst_mult_3_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_81 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[21]),
	.datac(!din_a[19]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_314 ),
	.cout(Xd_0__inst_mult_2_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_319 ),
	.cout(Xd_0__inst_mult_2_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_80 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[13]),
	.datac(!din_a[11]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_309 ),
	.cout(Xd_0__inst_mult_1_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_314 ),
	.cout(Xd_0__inst_mult_1_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_82 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[5]),
	.datac(!din_a[3]),
	.datad(!din_b[6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_319 ),
	.cout(Xd_0__inst_mult_0_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_324 ),
	.cout(Xd_0__inst_mult_0_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_83 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[253]),
	.datac(!din_a[252]),
	.datad(!din_b[254]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_324 ),
	.cout(Xd_0__inst_mult_31_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_82 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[237]),
	.datac(!din_a[236]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_319 ),
	.cout(Xd_0__inst_mult_29_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_83 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[229]),
	.datac(!din_a[228]),
	.datad(!din_b[230]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_324 ),
	.cout(Xd_0__inst_mult_28_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_82 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[221]),
	.datac(!din_a[220]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_319 ),
	.cout(Xd_0__inst_mult_27_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_81 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[117]),
	.datac(!din_a[116]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_313 ),
	.cout(Xd_0__inst_mult_14_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_82 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[109]),
	.datac(!din_a[108]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_318 ),
	.cout(Xd_0__inst_mult_13_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_81 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[101]),
	.datac(!din_a[100]),
	.datad(!din_b[102]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_313 ),
	.cout(Xd_0__inst_mult_12_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_82 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[93]),
	.datac(!din_a[92]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_318 ),
	.cout(Xd_0__inst_mult_11_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_82 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[85]),
	.datac(!din_a[84]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_318 ),
	.cout(Xd_0__inst_mult_10_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_81 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[77]),
	.datac(!din_a[76]),
	.datad(!din_b[78]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_313 ),
	.cout(Xd_0__inst_mult_9_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_82 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[69]),
	.datac(!din_a[68]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_318 ),
	.cout(Xd_0__inst_mult_8_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_81 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[61]),
	.datac(!din_a[60]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_313 ),
	.cout(Xd_0__inst_mult_7_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_82 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[53]),
	.datac(!din_a[52]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_318 ),
	.cout(Xd_0__inst_mult_6_319 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_81 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[45]),
	.datac(!din_a[44]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_309 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_313 ),
	.cout(Xd_0__inst_mult_5_314 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_83 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(!din_a[36]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_324 ),
	.cout(Xd_0__inst_mult_4_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_82 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[29]),
	.datac(!din_a[28]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_319 ),
	.cout(Xd_0__inst_mult_3_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_83 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[21]),
	.datac(!din_a[20]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_324 ),
	.cout(Xd_0__inst_mult_2_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_82 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[13]),
	.datac(!din_a[12]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_319 ),
	.cout(Xd_0__inst_mult_1_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_318 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_318 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_318 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_318 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_82 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_314 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_318 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_83 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_324 ),
	.cout(),
	.shareout());

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [16]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [17]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [18]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [19]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign [31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign [27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_31_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [31]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign [29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_27_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [27]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign [25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_23_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [23]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_19_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [19]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_30_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [30]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_28_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [28]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_29_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [29]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_31_ (
	.clk(clk),
	.d(Xd_0__inst_i21_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [31]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_26_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [26]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_24_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [24]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_25_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [25]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_27_ (
	.clk(clk),
	.d(Xd_0__inst_i21_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [27]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_22_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [22]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_20_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [20]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_21_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [21]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_23_ (
	.clk(clk),
	.d(Xd_0__inst_i21_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [23]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_18_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [18]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_16_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [16]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_17_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [17]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_19_ (
	.clk(clk),
	.d(Xd_0__inst_i21_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [19]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_15_ (
	.clk(clk),
	.d(Xd_0__inst_i21_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_11_ (
	.clk(clk),
	.d(Xd_0__inst_i21_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_7_ (
	.clk(clk),
	.d(Xd_0__inst_i21_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_3_ (
	.clk(clk),
	.d(Xd_0__inst_i21_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_113 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_109 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_118 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_114 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_123 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_119 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_133 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_129 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_138 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_134 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_30_ (
	.clk(clk),
	.d(Xd_0__inst_i21_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [30]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_28_ (
	.clk(clk),
	.d(Xd_0__inst_i21_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [28]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_29_ (
	.clk(clk),
	.d(Xd_0__inst_i21_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [29]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_26_ (
	.clk(clk),
	.d(Xd_0__inst_i21_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [26]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_24_ (
	.clk(clk),
	.d(Xd_0__inst_i21_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [24]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_25_ (
	.clk(clk),
	.d(Xd_0__inst_i21_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [25]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_22_ (
	.clk(clk),
	.d(Xd_0__inst_i21_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [22]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_20_ (
	.clk(clk),
	.d(Xd_0__inst_i21_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [20]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_21_ (
	.clk(clk),
	.d(Xd_0__inst_i21_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [21]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_18_ (
	.clk(clk),
	.d(Xd_0__inst_i21_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [18]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_16_ (
	.clk(clk),
	.d(Xd_0__inst_i21_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [16]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_17_ (
	.clk(clk),
	.d(Xd_0__inst_i21_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [17]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_14_ (
	.clk(clk),
	.d(Xd_0__inst_i21_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_12_ (
	.clk(clk),
	.d(Xd_0__inst_i21_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_13_ (
	.clk(clk),
	.d(Xd_0__inst_i21_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_10_ (
	.clk(clk),
	.d(Xd_0__inst_i21_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_143 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_8_ (
	.clk(clk),
	.d(Xd_0__inst_i21_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_9_ (
	.clk(clk),
	.d(Xd_0__inst_i21_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_6_ (
	.clk(clk),
	.d(Xd_0__inst_i21_131_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_4_ (
	.clk(clk),
	.d(Xd_0__inst_i21_136_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_5_ (
	.clk(clk),
	.d(Xd_0__inst_i21_141_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_2_ (
	.clk(clk),
	.d(Xd_0__inst_i21_146_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_0_ (
	.clk(clk),
	.d(Xd_0__inst_i21_151_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_1_ (
	.clk(clk),
	.d(Xd_0__inst_i21_156_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_139 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_153 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_158 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_149 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_154 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_154 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_154 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_178 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_183 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_154 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_159 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_193 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_164 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_198 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_203 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_174 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_179 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_213 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_189 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_218 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_223 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_194 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_199 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_233 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_209 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_14 (
	.clk(clk),
	.d(din_a[254]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_15 (
	.clk(clk),
	.d(din_b[251]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_14 (
	.clk(clk),
	.d(din_a[246]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_15 (
	.clk(clk),
	.d(din_b[243]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_14 (
	.clk(clk),
	.d(din_a[238]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_15 (
	.clk(clk),
	.d(din_b[235]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_14 (
	.clk(clk),
	.d(din_a[230]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_15 (
	.clk(clk),
	.d(din_b[227]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_14 (
	.clk(clk),
	.d(din_a[222]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_15 (
	.clk(clk),
	.d(din_b[219]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_14 (
	.clk(clk),
	.d(din_a[214]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_15 (
	.clk(clk),
	.d(din_b[211]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_14 (
	.clk(clk),
	.d(din_a[206]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_15 (
	.clk(clk),
	.d(din_b[203]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_14 (
	.clk(clk),
	.d(din_a[198]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_15 (
	.clk(clk),
	.d(din_b[195]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_14 (
	.clk(clk),
	.d(din_a[190]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_15 (
	.clk(clk),
	.d(din_b[187]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_14 (
	.clk(clk),
	.d(din_a[182]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_15 (
	.clk(clk),
	.d(din_b[179]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_14 (
	.clk(clk),
	.d(din_a[174]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_15 (
	.clk(clk),
	.d(din_b[171]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_14 (
	.clk(clk),
	.d(din_a[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_15 (
	.clk(clk),
	.d(din_b[163]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_14 (
	.clk(clk),
	.d(din_a[158]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_15 (
	.clk(clk),
	.d(din_b[155]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_14 (
	.clk(clk),
	.d(din_a[150]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_15 (
	.clk(clk),
	.d(din_b[147]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_14 (
	.clk(clk),
	.d(din_a[142]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_15 (
	.clk(clk),
	.d(din_b[139]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_14 (
	.clk(clk),
	.d(din_a[134]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_15 (
	.clk(clk),
	.d(din_b[131]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_14 (
	.clk(clk),
	.d(din_a[126]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_15 (
	.clk(clk),
	.d(din_b[123]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_14 (
	.clk(clk),
	.d(din_a[118]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_15 (
	.clk(clk),
	.d(din_b[115]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_14 (
	.clk(clk),
	.d(din_a[110]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_15 (
	.clk(clk),
	.d(din_b[107]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_14 (
	.clk(clk),
	.d(din_a[102]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_15 (
	.clk(clk),
	.d(din_b[99]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_14 (
	.clk(clk),
	.d(din_a[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_15 (
	.clk(clk),
	.d(din_b[91]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_14 (
	.clk(clk),
	.d(din_a[86]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_15 (
	.clk(clk),
	.d(din_b[83]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_14 (
	.clk(clk),
	.d(din_a[78]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_15 (
	.clk(clk),
	.d(din_b[75]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_14 (
	.clk(clk),
	.d(din_a[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_15 (
	.clk(clk),
	.d(din_b[67]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_14 (
	.clk(clk),
	.d(din_a[62]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_15 (
	.clk(clk),
	.d(din_b[59]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_14 (
	.clk(clk),
	.d(din_a[54]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_15 (
	.clk(clk),
	.d(din_b[51]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_238 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_243 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_14 (
	.clk(clk),
	.d(din_a[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_15 (
	.clk(clk),
	.d(din_b[43]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_14 (
	.clk(clk),
	.d(din_a[38]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_15 (
	.clk(clk),
	.d(din_b[35]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_14 (
	.clk(clk),
	.d(din_a[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_15 (
	.clk(clk),
	.d(din_b[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_14 (
	.clk(clk),
	.d(din_a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_15 (
	.clk(clk),
	.d(din_b[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_14 (
	.clk(clk),
	.d(din_a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_15 (
	.clk(clk),
	.d(din_b[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_14 (
	.clk(clk),
	.d(din_a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_15 (
	.clk(clk),
	.d(din_b[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_263 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_263 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_263 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_263 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_263 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_253 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_23_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_263 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_258 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_28_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_21_q ));

assign dout[0] = Xd_0__inst_inst_inst_inst_dout [0];

assign dout[1] = Xd_0__inst_inst_inst_inst_dout [1];

assign dout[2] = Xd_0__inst_inst_inst_inst_dout [2];

assign dout[3] = Xd_0__inst_inst_inst_inst_dout [3];

assign dout[4] = Xd_0__inst_inst_inst_inst_dout [4];

assign dout[5] = Xd_0__inst_inst_inst_inst_dout [5];

assign dout[6] = Xd_0__inst_inst_inst_inst_dout [6];

assign dout[7] = Xd_0__inst_inst_inst_inst_dout [7];

assign dout[8] = Xd_0__inst_inst_inst_inst_dout [8];

assign dout[9] = Xd_0__inst_inst_inst_inst_dout [9];

assign dout[10] = Xd_0__inst_inst_inst_inst_dout [10];

assign dout[11] = Xd_0__inst_inst_inst_inst_dout [11];

assign dout[12] = Xd_0__inst_inst_inst_inst_dout [12];

assign dout[13] = Xd_0__inst_inst_inst_inst_dout [13];

assign dout[14] = Xd_0__inst_inst_inst_inst_dout [14];

assign dout[15] = Xd_0__inst_inst_inst_inst_dout [15];

assign dout[16] = Xd_0__inst_inst_inst_inst_dout [16];

assign dout[17] = Xd_0__inst_inst_inst_inst_dout [17];

assign dout[18] = Xd_0__inst_inst_inst_inst_dout [18];

assign dout[19] = Xd_0__inst_inst_inst_inst_dout [19];

endmodule
